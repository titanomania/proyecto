library IEEE;
use IEEE.std_logic_1164.all;

entity Mux256a18Bits is
    port (
        d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15,
        d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31,
        d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47,
        d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63,
        d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79,
        d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95,
        d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111,
        d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127,
        d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143,
        d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159,
        d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175,
        d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191,
        d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207,
        d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223,
        d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239,
        d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255: in std_logic_vector(7 downto 0);
        S: in std_logic_vector(7 downto 0);
        r: out std_logic_vector(7 downto 0)
    );
end Mux256a18Bits;

architecture Ar_Mux256a18Bits of Mux256a18Bits is
    
    component Mux256a1 is
        port (
            d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15,
            d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31,
            d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47,
            d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63,
            d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79,
            d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95,
            d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111,
            d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127,
            d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143,
            d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159,
            d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175,
            d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191,
            d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207,
            d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223,
            d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239,
            d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255: in std_logic;
            S: in std_logic_vector (7 downto 0);
            r: out std_logic
        );
    end component;

    begin
        Mux256a1_0: Mux256a1 port map (d0(0), d1(0), d2(0), d3(0), d4(0), d5(0), d6(0), d7(0),
            d8(0), d9(0), d10(0), d11(0), d12(0), d13(0), d14(0), d15(0),
            d16(0), d17(0), d18(0), d19(0), d20(0), d21(0), d22(0), d23(0),
            d24(0), d25(0), d26(0), d27(0), d28(0), d29(0), d30(0), d31(0),
            d32(0), d33(0), d34(0), d35(0), d36(0), d37(0), d38(0), d39(0),
            d40(0), d41(0), d42(0), d43(0), d44(0), d45(0), d46(0), d47(0),
            d48(0), d49(0), d50(0), d51(0), d52(0), d53(0), d54(0), d55(0),
            d56(0), d57(0), d58(0), d59(0), d60(0), d61(0), d62(0), d63(0),
            d64(0), d65(0), d66(0), d67(0), d68(0), d69(0), d70(0), d71(0),
            d72(0), d73(0), d74(0), d75(0), d76(0), d77(0), d78(0), d79(0),
            d80(0), d81(0), d82(0), d83(0), d84(0), d85(0), d86(0), d87(0),
            d88(0), d89(0), d90(0), d91(0), d92(0), d93(0), d94(0), d95(0),
            d96(0), d97(0), d98(0), d99(0), d100(0), d101(0), d102(0), d103(0),
            d104(0), d105(0), d106(0), d107(0), d108(0), d109(0), d110(0), d111(0),
            d112(0), d113(0), d114(0), d115(0), d116(0), d117(0), d118(0), d119(0),
            d120(0), d121(0), d122(0), d123(0), d124(0), d125(0), d126(0), d127(0),
            d128(0), d129(0), d130(0), d131(0), d132(0), d133(0), d134(0), d135(0),
            d136(0), d137(0), d138(0), d139(0), d140(0), d141(0), d142(0), d143(0),
            d144(0), d145(0), d146(0), d147(0), d148(0), d149(0), d150(0), d151(0),
            d152(0), d153(0), d154(0), d155(0), d156(0), d157(0), d158(0), d159(0),
            d160(0), d161(0), d162(0), d163(0), d164(0), d165(0), d166(0), d167(0),
            d168(0), d169(0), d170(0), d171(0), d172(0), d173(0), d174(0), d175(0),
            d176(0), d177(0), d178(0), d179(0), d180(0), d181(0), d182(0), d183(0),
            d184(0), d185(0), d186(0), d187(0), d188(0), d189(0), d190(0), d191(0),
            d192(0), d193(0), d194(0), d195(0), d196(0), d197(0), d198(0), d199(0),
            d200(0), d201(0), d202(0), d203(0), d204(0), d205(0), d206(0), d207(0),
            d208(0), d209(0), d210(0), d211(0), d212(0), d213(0), d214(0), d215(0),
            d216(0), d217(0), d218(0), d219(0), d220(0), d221(0), d222(0), d223(0),
            d224(0), d225(0), d226(0), d227(0), d228(0), d229(0), d230(0), d231(0),
            d232(0), d233(0), d234(0), d235(0), d236(0), d237(0), d238(0), d239(0),
            d240(0), d241(0), d242(0), d243(0), d244(0), d245(0), d246(0), d247(0),
            d248(0), d249(0), d250(0), d251(0), d252(0), d253(0), d254(0), d255(0),
            S,
            r (0)
        );

        Mux256a1_1: Mux256a1 port map (d0(1), d1(1), d2(1), d3(1), d4(1), d5(1), d6(1), d7(1),
            d8(1), d9(1), d10(1), d11(1), d12(1), d13(1), d14(1), d15(1),
            d16(1), d17(1), d18(1), d19(1), d20(1), d21(1), d22(1), d23(1),
            d24(1), d25(1), d26(1), d27(1), d28(1), d29(1), d30(1), d31(1),
            d32(1), d33(1), d34(1), d35(1), d36(1), d37(1), d38(1), d39(1),
            d40(1), d41(1), d42(1), d43(1), d44(1), d45(1), d46(1), d47(1),
            d48(1), d49(1), d50(1), d51(1), d52(1), d53(1), d54(1), d55(1),
            d56(1), d57(1), d58(1), d59(1), d60(1), d61(1), d62(1), d63(1),
            d64(1), d65(1), d66(1), d67(1), d68(1), d69(1), d70(1), d71(1),
            d72(1), d73(1), d74(1), d75(1), d76(1), d77(1), d78(1), d79(1),
            d80(1), d81(1), d82(1), d83(1), d84(1), d85(1), d86(1), d87(1),
            d88(1), d89(1), d90(1), d91(1), d92(1), d93(1), d94(1), d95(1),
            d96(1), d97(1), d98(1), d99(1), d100(1), d101(1), d102(1), d103(1),
            d104(1), d105(1), d106(1), d107(1), d108(1), d109(1), d110(1), d111(1),
            d112(1), d113(1), d114(1), d115(1), d116(1), d117(1), d118(1), d119(1),
            d120(1), d121(1), d122(1), d123(1), d124(1), d125(1), d126(1), d127(1),
            d128(1), d129(1), d130(1), d131(1), d132(1), d133(1), d134(1), d135(1),
            d136(1), d137(1), d138(1), d139(1), d140(1), d141(1), d142(1), d143(1),
            d144(1), d145(1), d146(1), d147(1), d148(1), d149(1), d150(1), d151(1),
            d152(1), d153(1), d154(1), d155(1), d156(1), d157(1), d158(1), d159(1),
            d160(1), d161(1), d162(1), d163(1), d164(1), d165(1), d166(1), d167(1),
            d168(1), d169(1), d170(1), d171(1), d172(1), d173(1), d174(1), d175(1),
            d176(1), d177(1), d178(1), d179(1), d180(1), d181(1), d182(1), d183(1),
            d184(1), d185(1), d186(1), d187(1), d188(1), d189(1), d190(1), d191(1),
            d192(1), d193(1), d194(1), d195(1), d196(1), d197(1), d198(1), d199(1),
            d200(1), d201(1), d202(1), d203(1), d204(1), d205(1), d206(1), d207(1),
            d208(1), d209(1), d210(1), d211(1), d212(1), d213(1), d214(1), d215(1),
            d216(1), d217(1), d218(1), d219(1), d220(1), d221(1), d222(1), d223(1),
            d224(1), d225(1), d226(1), d227(1), d228(1), d229(1), d230(1), d231(1),
            d232(1), d233(1), d234(1), d235(1), d236(1), d237(1), d238(1), d239(1),
            d240(1), d241(1), d242(1), d243(1), d244(1), d245(1), d246(1), d247(1),
            d248(1), d249(1), d250(1), d251(1), d252(1), d253(1), d254(1), d255(1),
            S,
            r (1)
        );

        Mux256a1_2: Mux256a1 port map (d0(2), d1(2), d2(2), d3(2), d4(2), d5(2), d6(2), d7(2),
            d8(2), d9(2), d10(2), d11(2), d12(2), d13(2), d14(2), d15(2),
            d16(2), d17(2), d18(2), d19(2), d20(2), d21(2), d22(2), d23(2),
            d24(2), d25(2), d26(2), d27(2), d28(2), d29(2), d30(2), d31(2),
            d32(2), d33(2), d34(2), d35(2), d36(2), d37(2), d38(2), d39(2),
            d40(2), d41(2), d42(2), d43(2), d44(2), d45(2), d46(2), d47(2),
            d48(2), d49(2), d50(2), d51(2), d52(2), d53(2), d54(2), d55(2),
            d56(2), d57(2), d58(2), d59(2), d60(2), d61(2), d62(2), d63(2),
            d64(2), d65(2), d66(2), d67(2), d68(2), d69(2), d70(2), d71(2),
            d72(2), d73(2), d74(2), d75(2), d76(2), d77(2), d78(2), d79(2),
            d80(2), d81(2), d82(2), d83(2), d84(2), d85(2), d86(2), d87(2),
            d88(2), d89(2), d90(2), d91(2), d92(2), d93(2), d94(2), d95(2),
            d96(2), d97(2), d98(2), d99(2), d100(2), d101(2), d102(2), d103(2),
            d104(2), d105(2), d106(2), d107(2), d108(2), d109(2), d110(2), d111(2),
            d112(2), d113(2), d114(2), d115(2), d116(2), d117(2), d118(2), d119(2),
            d120(2), d121(2), d122(2), d123(2), d124(2), d125(2), d126(2), d127(2),
            d128(2), d129(2), d130(2), d131(2), d132(2), d133(2), d134(2), d135(2),
            d136(2), d137(2), d138(2), d139(2), d140(2), d141(2), d142(2), d143(2),
            d144(2), d145(2), d146(2), d147(2), d148(2), d149(2), d150(2), d151(2),
            d152(2), d153(2), d154(2), d155(2), d156(2), d157(2), d158(2), d159(2),
            d160(2), d161(2), d162(2), d163(2), d164(2), d165(2), d166(2), d167(2),
            d168(2), d169(2), d170(2), d171(2), d172(2), d173(2), d174(2), d175(2),
            d176(2), d177(2), d178(2), d179(2), d180(2), d181(2), d182(2), d183(2),
            d184(2), d185(2), d186(2), d187(2), d188(2), d189(2), d190(2), d191(2),
            d192(2), d193(2), d194(2), d195(2), d196(2), d197(2), d198(2), d199(2),
            d200(2), d201(2), d202(2), d203(2), d204(2), d205(2), d206(2), d207(2),
            d208(2), d209(2), d210(2), d211(2), d212(2), d213(2), d214(2), d215(2),
            d216(2), d217(2), d218(2), d219(2), d220(2), d221(2), d222(2), d223(2),
            d224(2), d225(2), d226(2), d227(2), d228(2), d229(2), d230(2), d231(2),
            d232(2), d233(2), d234(2), d235(2), d236(2), d237(2), d238(2), d239(2),
            d240(2), d241(2), d242(2), d243(2), d244(2), d245(2), d246(2), d247(2),
            d248(2), d249(2), d250(2), d251(2), d252(2), d253(2), d254(2), d255(2),
            S,
            r (2)
        );

        Mux256a1_3: Mux256a1 port map (d0(3), d1(3), d2(3), d3(3), d4(3), d5(3), d6(3), d7(3),
            d8(3), d9(3), d10(3), d11(3), d12(3), d13(3), d14(3), d15(3),
            d16(3), d17(3), d18(3), d19(3), d20(3), d21(3), d22(3), d23(3),
            d24(3), d25(3), d26(3), d27(3), d28(3), d29(3), d30(3), d31(3),
            d32(3), d33(3), d34(3), d35(3), d36(3), d37(3), d38(3), d39(3),
            d40(3), d41(3), d42(3), d43(3), d44(3), d45(3), d46(3), d47(3),
            d48(3), d49(3), d50(3), d51(3), d52(3), d53(3), d54(3), d55(3),
            d56(3), d57(3), d58(3), d59(3), d60(3), d61(3), d62(3), d63(3),
            d64(3), d65(3), d66(3), d67(3), d68(3), d69(3), d70(3), d71(3),
            d72(3), d73(3), d74(3), d75(3), d76(3), d77(3), d78(3), d79(3),
            d80(3), d81(3), d82(3), d83(3), d84(3), d85(3), d86(3), d87(3),
            d88(3), d89(3), d90(3), d91(3), d92(3), d93(3), d94(3), d95(3),
            d96(3), d97(3), d98(3), d99(3), d100(3), d101(3), d102(3), d103(3),
            d104(3), d105(3), d106(3), d107(3), d108(3), d109(3), d110(3), d111(3),
            d112(3), d113(3), d114(3), d115(3), d116(3), d117(3), d118(3), d119(3),
            d120(3), d121(3), d122(3), d123(3), d124(3), d125(3), d126(3), d127(3),
            d128(3), d129(3), d130(3), d131(3), d132(3), d133(3), d134(3), d135(3),
            d136(3), d137(3), d138(3), d139(3), d140(3), d141(3), d142(3), d143(3),
            d144(3), d145(3), d146(3), d147(3), d148(3), d149(3), d150(3), d151(3),
            d152(3), d153(3), d154(3), d155(3), d156(3), d157(3), d158(3), d159(3),
            d160(3), d161(3), d162(3), d163(3), d164(3), d165(3), d166(3), d167(3),
            d168(3), d169(3), d170(3), d171(3), d172(3), d173(3), d174(3), d175(3),
            d176(3), d177(3), d178(3), d179(3), d180(3), d181(3), d182(3), d183(3),
            d184(3), d185(3), d186(3), d187(3), d188(3), d189(3), d190(3), d191(3),
            d192(3), d193(3), d194(3), d195(3), d196(3), d197(3), d198(3), d199(3),
            d200(3), d201(3), d202(3), d203(3), d204(3), d205(3), d206(3), d207(3),
            d208(3), d209(3), d210(3), d211(3), d212(3), d213(3), d214(3), d215(3),
            d216(3), d217(3), d218(3), d219(3), d220(3), d221(3), d222(3), d223(3),
            d224(3), d225(3), d226(3), d227(3), d228(3), d229(3), d230(3), d231(3),
            d232(3), d233(3), d234(3), d235(3), d236(3), d237(3), d238(3), d239(3),
            d240(3), d241(3), d242(3), d243(3), d244(3), d245(3), d246(3), d247(3),
            d248(3), d249(3), d250(3), d251(3), d252(3), d253(3), d254(3), d255(3),
            S,
            r (3)
        );

        
        Mux256a1_4: Mux256a1 port map (d0(4), d1(4), d2(4), d3(4), d4(4), d5(4), d6(4), d7(4),
            d8(4), d9(4), d10(4), d11(4), d12(4), d13(4), d14(4), d15(4),
            d16(4), d17(4), d18(4), d19(4), d20(4), d21(4), d22(4), d23(4),
            d24(4), d25(4), d26(4), d27(4), d28(4), d29(4), d30(4), d31(4),
            d32(4), d33(4), d34(4), d35(4), d36(4), d37(4), d38(4), d39(4),
            d40(4), d41(4), d42(4), d43(4), d44(4), d45(4), d46(4), d47(4),
            d48(4), d49(4), d50(4), d51(4), d52(4), d53(4), d54(4), d55(4),
            d56(4), d57(4), d58(4), d59(4), d60(4), d61(4), d62(4), d63(4),
            d64(4), d65(4), d66(4), d67(4), d68(4), d69(4), d70(4), d71(4),
            d72(4), d73(4), d74(4), d75(4), d76(4), d77(4), d78(4), d79(4),
            d80(4), d81(4), d82(4), d83(4), d84(4), d85(4), d86(4), d87(4),
            d88(4), d89(4), d90(4), d91(4), d92(4), d93(4), d94(4), d95(4),
            d96(4), d97(4), d98(4), d99(4), d100(4), d101(4), d102(4), d103(4),
            d104(4), d105(4), d106(4), d107(4), d108(4), d109(4), d110(4), d111(4),
            d112(4), d113(4), d114(4), d115(4), d116(4), d117(4), d118(4), d119(4),
            d120(4), d121(4), d122(4), d123(4), d124(4), d125(4), d126(4), d127(4),
            d128(4), d129(4), d130(4), d131(4), d132(4), d133(4), d134(4), d135(4),
            d136(4), d137(4), d138(4), d139(4), d140(4), d141(4), d142(4), d143(4),
            d144(4), d145(4), d146(4), d147(4), d148(4), d149(4), d150(4), d151(4),
            d152(4), d153(4), d154(4), d155(4), d156(4), d157(4), d158(4), d159(4),
            d160(4), d161(4), d162(4), d163(4), d164(4), d165(4), d166(4), d167(4),
            d168(4), d169(4), d170(4), d171(4), d172(4), d173(4), d174(4), d175(4),
            d176(4), d177(4), d178(4), d179(4), d180(4), d181(4), d182(4), d183(4),
            d184(4), d185(4), d186(4), d187(4), d188(4), d189(4), d190(4), d191(4),
            d192(4), d193(4), d194(4), d195(4), d196(4), d197(4), d198(4), d199(4),
            d200(4), d201(4), d202(4), d203(4), d204(4), d205(4), d206(4), d207(4),
            d208(4), d209(4), d210(4), d211(4), d212(4), d213(4), d214(4), d215(4),
            d216(4), d217(4), d218(4), d219(4), d220(4), d221(4), d222(4), d223(4),
            d224(4), d225(4), d226(4), d227(4), d228(4), d229(4), d230(4), d231(4),
            d232(4), d233(4), d234(4), d235(4), d236(4), d237(4), d238(4), d239(4),
            d240(4), d241(4), d242(4), d243(4), d244(4), d245(4), d246(4), d247(4),
            d248(4), d249(4), d250(4), d251(4), d252(4), d253(4), d254(4), d255(4),
            S,
            r (4)
        );

        Mux256a1_5: Mux256a1 port map (d0(5), d1(5), d2(5), d3(5), d4(5), d5(5), d6(5), d7(5),
            d8(5), d9(5), d10(5), d11(5), d12(5), d13(5), d14(5), d15(5),
            d16(5), d17(5), d18(5), d19(5), d20(5), d21(5), d22(5), d23(5),
            d24(5), d25(5), d26(5), d27(5), d28(5), d29(5), d30(5), d31(5),
            d32(5), d33(5), d34(5), d35(5), d36(5), d37(5), d38(5), d39(5),
            d40(5), d41(5), d42(5), d43(5), d44(5), d45(5), d46(5), d47(5),
            d48(5), d49(5), d50(5), d51(5), d52(5), d53(5), d54(5), d55(5),
            d56(5), d57(5), d58(5), d59(5), d60(5), d61(5), d62(5), d63(5),
            d64(5), d65(5), d66(5), d67(5), d68(5), d69(5), d70(5), d71(5),
            d72(5), d73(5), d74(5), d75(5), d76(5), d77(5), d78(5), d79(5),
            d80(5), d81(5), d82(5), d83(5), d84(5), d85(5), d86(5), d87(5),
            d88(5), d89(5), d90(5), d91(5), d92(5), d93(5), d94(5), d95(5),
            d96(5), d97(5), d98(5), d99(5), d100(5), d101(5), d102(5), d103(5),
            d104(5), d105(5), d106(5), d107(5), d108(5), d109(5), d110(5), d111(5),
            d112(5), d113(5), d114(5), d115(5), d116(5), d117(5), d118(5), d119(5),
            d120(5), d121(5), d122(5), d123(5), d124(5), d125(5), d126(5), d127(5),
            d128(5), d129(5), d130(5), d131(5), d132(5), d133(5), d134(5), d135(5),
            d136(5), d137(5), d138(5), d139(5), d140(5), d141(5), d142(5), d143(5),
            d144(5), d145(5), d146(5), d147(5), d148(5), d149(5), d150(5), d151(5),
            d152(5), d153(5), d154(5), d155(5), d156(5), d157(5), d158(5), d159(5),
            d160(5), d161(5), d162(5), d163(5), d164(5), d165(5), d166(5), d167(5),
            d168(5), d169(5), d170(5), d171(5), d172(5), d173(5), d174(5), d175(5),
            d176(5), d177(5), d178(5), d179(5), d180(5), d181(5), d182(5), d183(5),
            d184(5), d185(5), d186(5), d187(5), d188(5), d189(5), d190(5), d191(5),
            d192(5), d193(5), d194(5), d195(5), d196(5), d197(5), d198(5), d199(5),
            d200(5), d201(5), d202(5), d203(5), d204(5), d205(5), d206(5), d207(5),
            d208(5), d209(5), d210(5), d211(5), d212(5), d213(5), d214(5), d215(5),
            d216(5), d217(5), d218(5), d219(5), d220(5), d221(5), d222(5), d223(5),
            d224(5), d225(5), d226(5), d227(5), d228(5), d229(5), d230(5), d231(5),
            d232(5), d233(5), d234(5), d235(5), d236(5), d237(5), d238(5), d239(5),
            d240(5), d241(5), d242(5), d243(5), d244(5), d245(5), d246(5), d247(5),
            d248(5), d249(5), d250(5), d251(5), d252(5), d253(5), d254(5), d255(5),
            S,
            r (5)
        );

        Mux256a1_6: Mux256a1 port map (d0(6), d1(6), d2(6), d3(6), d4(6), d5(6), d6(6), d7(6),
            d8(6), d9(6), d10(6), d11(6), d12(6), d13(6), d14(6), d15(6),
            d16(6), d17(6), d18(6), d19(6), d20(6), d21(6), d22(6), d23(6),
            d24(6), d25(6), d26(6), d27(6), d28(6), d29(6), d30(6), d31(6),
            d32(6), d33(6), d34(6), d35(6), d36(6), d37(6), d38(6), d39(6),
            d40(6), d41(6), d42(6), d43(6), d44(6), d45(6), d46(6), d47(6),
            d48(6), d49(6), d50(6), d51(6), d52(6), d53(6), d54(6), d55(6),
            d56(6), d57(6), d58(6), d59(6), d60(6), d61(6), d62(6), d63(6),
            d64(6), d65(6), d66(6), d67(6), d68(6), d69(6), d70(6), d71(6),
            d72(6), d73(6), d74(6), d75(6), d76(6), d77(6), d78(6), d79(6),
            d80(6), d81(6), d82(6), d83(6), d84(6), d85(6), d86(6), d87(6),
            d88(6), d89(6), d90(6), d91(6), d92(6), d93(6), d94(6), d95(6),
            d96(6), d97(6), d98(6), d99(6), d100(6), d101(6), d102(6), d103(6),
            d104(6), d105(6), d106(6), d107(6), d108(6), d109(6), d110(6), d111(6),
            d112(6), d113(6), d114(6), d115(6), d116(6), d117(6), d118(6), d119(6),
            d120(6), d121(6), d122(6), d123(6), d124(6), d125(6), d126(6), d127(6),
            d128(6), d129(6), d130(6), d131(6), d132(6), d133(6), d134(6), d135(6),
            d136(6), d137(6), d138(6), d139(6), d140(6), d141(6), d142(6), d143(6),
            d144(6), d145(6), d146(6), d147(6), d148(6), d149(6), d150(6), d151(6),
            d152(6), d153(6), d154(6), d155(6), d156(6), d157(6), d158(6), d159(6),
            d160(6), d161(6), d162(6), d163(6), d164(6), d165(6), d166(6), d167(6),
            d168(6), d169(6), d170(6), d171(6), d172(6), d173(6), d174(6), d175(6),
            d176(6), d177(6), d178(6), d179(6), d180(6), d181(6), d182(6), d183(6),
            d184(6), d185(6), d186(6), d187(6), d188(6), d189(6), d190(6), d191(6),
            d192(6), d193(6), d194(6), d195(6), d196(6), d197(6), d198(6), d199(6),
            d200(6), d201(6), d202(6), d203(6), d204(6), d205(6), d206(6), d207(6),
            d208(6), d209(6), d210(6), d211(6), d212(6), d213(6), d214(6), d215(6),
            d216(6), d217(6), d218(6), d219(6), d220(6), d221(6), d222(6), d223(6),
            d224(6), d225(6), d226(6), d227(6), d228(6), d229(6), d230(6), d231(6),
            d232(6), d233(6), d234(6), d235(6), d236(6), d237(6), d238(6), d239(6),
            d240(6), d241(6), d242(6), d243(6), d244(6), d245(6), d246(6), d247(6),
            d248(6), d249(6), d250(6), d251(6), d252(6), d253(6), d254(6), d255(6),
            S,
            r (6)
        );

        Mux256a1_7: Mux256a1 port map (d0(7), d1(7), d2(7), d3(7), d4(7), d5(7), d6(7), d7(7),
            d8(7), d9(7), d10(7), d11(7), d12(7), d13(7), d14(7), d15(7),
            d16(7), d17(7), d18(7), d19(7), d20(7), d21(7), d22(7), d23(7),
            d24(7), d25(7), d26(7), d27(7), d28(7), d29(7), d30(7), d31(7),
            d32(7), d33(7), d34(7), d35(7), d36(7), d37(7), d38(7), d39(7),
            d40(7), d41(7), d42(7), d43(7), d44(7), d45(7), d46(7), d47(7),
            d48(7), d49(7), d50(7), d51(7), d52(7), d53(7), d54(7), d55(7),
            d56(7), d57(7), d58(7), d59(7), d60(7), d61(7), d62(7), d63(7),
            d64(7), d65(7), d66(7), d67(7), d68(7), d69(7), d70(7), d71(7),
            d72(7), d73(7), d74(7), d75(7), d76(7), d77(7), d78(7), d79(7),
            d80(7), d81(7), d82(7), d83(7), d84(7), d85(7), d86(7), d87(7),
            d88(7), d89(7), d90(7), d91(7), d92(7), d93(7), d94(7), d95(7),
            d96(7), d97(7), d98(7), d99(7), d100(7), d101(7), d102(7), d103(7),
            d104(7), d105(7), d106(7), d107(7), d108(7), d109(7), d110(7), d111(7),
            d112(7), d113(7), d114(7), d115(7), d116(7), d117(7), d118(7), d119(7),
            d120(7), d121(7), d122(7), d123(7), d124(7), d125(7), d126(7), d127(7),
            d128(7), d129(7), d130(7), d131(7), d132(7), d133(7), d134(7), d135(7),
            d136(7), d137(7), d138(7), d139(7), d140(7), d141(7), d142(7), d143(7),
            d144(7), d145(7), d146(7), d147(7), d148(7), d149(7), d150(7), d151(7),
            d152(7), d153(7), d154(7), d155(7), d156(7), d157(7), d158(7), d159(7),
            d160(7), d161(7), d162(7), d163(7), d164(7), d165(7), d166(7), d167(7),
            d168(7), d169(7), d170(7), d171(7), d172(7), d173(7), d174(7), d175(7),
            d176(7), d177(7), d178(7), d179(7), d180(7), d181(7), d182(7), d183(7),
            d184(7), d185(7), d186(7), d187(7), d188(7), d189(7), d190(7), d191(7),
            d192(7), d193(7), d194(7), d195(7), d196(7), d197(7), d198(7), d199(7),
            d200(7), d201(7), d202(7), d203(7), d204(7), d205(7), d206(7), d207(7),
            d208(7), d209(7), d210(7), d211(7), d212(7), d213(7), d214(7), d215(7),
            d216(7), d217(7), d218(7), d219(7), d220(7), d221(7), d222(7), d223(7),
            d224(7), d225(7), d226(7), d227(7), d228(7), d229(7), d230(7), d231(7),
            d232(7), d233(7), d234(7), d235(7), d236(7), d237(7), d238(7), d239(7),
            d240(7), d241(7), d242(7), d243(7), d244(7), d245(7), d246(7), d247(7),
            d248(7), d249(7), d250(7), d251(7), d252(7), d253(7), d254(7), d255(7),
            S,
            r (7)
        );



    end architecture;