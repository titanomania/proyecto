library IEEE;
use IEEE.std_logic_1164.all;

entity Deco8a256 is
  port (
    S: in std_logic_vector(7 downto 0);
    d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15,
          d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31,
          d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47,
          d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63,
          d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79,
          d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95,
          d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111,
          d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127,
          d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143,
          d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159,
          d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175,
          d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191,
          d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207,
          d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223,
          d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239,
          d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255: out std_logic
  );
end Deco8a256;

architecture Ar_Deco8a256 of Deco8a256 is
begin

    d0   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d1   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d2   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d3   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d4   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d5   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d6   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d7   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d8   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d9   <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d10  <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d11  <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d12  <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d13  <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d14  <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d15  <= not(S(7)) and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d16  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d17  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d18  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d19  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d20  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d21  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d22  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d23  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d24  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d25  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d26  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d27  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d28  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d29  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d30  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d31  <= not(S(7)) and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and S(0);
    d32  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d33  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d34  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d35  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d36  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d37  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d38  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d39  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d40  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d41  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d42  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d43  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d44  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d45  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d46  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d47  <= not(S(7)) and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d48  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d49  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d50  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d51  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d52  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d53  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d54  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d55  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d56  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d57  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d58  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d59  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d60  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d61  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d62  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d63  <= not(S(7)) and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and S(0);
    d64  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d65  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d66  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d67  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d68  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d69  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d70  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d71  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d72  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d73  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d74  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d75  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d76  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d77  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d78  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d79  <= not(S(7)) and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d80  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d81  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d82  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d83  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d84  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d85  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d86  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d87  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d88  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d89  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d90  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d91  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d92  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d93  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d94  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d95  <= not(S(7)) and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and S(0);
    d96  <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d97  <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d98  <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d99  <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d100 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d101 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d102 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d103 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d104 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d105 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d106 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d107 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d108 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d109 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d110 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d111 <= not(S(7)) and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d112 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d113 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d114 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d115 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d116 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d117 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d118 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d119 <= not(S(7)) and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d120 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d121 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d122 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d123 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d124 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d125 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d126 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d127 <= not(S(7)) and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and S(0);
    d128 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d129 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d130 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d131 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d132 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d133 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d134 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d135 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d136 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d137 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d138 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d139 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d140 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d141 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d142 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d143 <= S(7)      and not(S(6)) and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d144 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d145 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d146 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d147 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d148 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d149 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d150 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d151 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d152 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d153 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d154 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d155 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d156 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d157 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d158 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d159 <= S(7)      and not(S(6)) and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and S(0);
    d160 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d161 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d162 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d163 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d164 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d165 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d166 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d167 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d168 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d169 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d170 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d171 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d172 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d173 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d174 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d175 <= S(7)      and not(S(6)) and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d176 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d177 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d178 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d179 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d180 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d181 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d182 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d183 <= S(7)      and not(S(6)) and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d184 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d185 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d186 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d187 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d188 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d189 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d190 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d191 <= S(7)      and not(S(6)) and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and S(0);
    d192 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d193 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d194 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d195 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d196 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d197 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d198 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d199 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d200 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d201 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d202 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d203 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d204 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d205 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d206 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d207 <= S(7)      and S(6)      and not(S(5)) and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d208 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d209 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d210 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d211 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d212 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d213 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d214 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d215 <= S(7)      and S(6)      and not(S(5)) and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d216 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d217 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d218 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d219 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d220 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d221 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d222 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d223 <= S(7)      and S(6)      and not(S(5)) and S(4)      and S(3)      and S(2)      and S(1)      and S(0);
    d224 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d225 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d226 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d227 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d228 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d229 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d230 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d231 <= S(7)      and S(6)      and S(5)      and not(S(4)) and not(S(3)) and S(2)      and S(1)      and S(0);
    d232 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d233 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d234 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d235 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and not(S(2)) and S(1)      and S(0);
    d236 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d237 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and not(S(1)) and S(0);
    d238 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and not(S(0));
    d239 <= S(7)      and S(6)      and S(5)      and not(S(4)) and S(3)      and S(2)      and S(1)      and S(0);
    d240 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and not(S(0));
    d241 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and not(S(1)) and S(0);
    d242 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and not(S(0));
    d243 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and not(S(2)) and S(1)      and S(0);
    d244 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and not(S(0));
    d245 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and not(S(1)) and S(0);
    d246 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and not(S(0));
    d247 <= S(7)      and S(6)      and S(5)      and S(4)      and not(S(3)) and S(2)      and S(1)      and S(0);
    d248 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and not(S(0));
    d249 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and not(S(1)) and S(0);
    d250 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and not(S(0));
    d251 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and not(S(2)) and S(1)      and S(0);
    d252 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and not(S(0));
    d253 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and not(S(1)) and S(0);
    d254 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and not(S(0));
    d255 <= S(7)      and S(6)      and S(5)      and S(4)      and S(3)      and S(2)      and S(1)      and S(0);




end Ar_Deco8a256;
