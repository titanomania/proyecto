library IEEE;
use IEEE.std_logic_1164.all;

entity Mux256a125Bits is
    port (
        d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15,
        d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31,
        d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47,
        d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63,
        d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79,
        d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95,
        d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111,
        d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127,
        d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143,
        d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159,
        d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175,
        d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191,
        d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207,
        d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223,
        d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239,
        d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255: in std_logic_vector(24 downto 0);
        S: in std_logic_vector(7 downto 0);
        r: out std_logic_vector(24 downto 0)
    );
end Mux256a125Bits;

architecture Ar_Mux256a125Bits of Mux256a125Bits is
    
    component Mux256a1 is
        port (
            d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15,
            d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31,
            d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47,
            d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63,
            d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79,
            d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95,
            d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111,
            d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127,
            d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143,
            d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159,
            d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175,
            d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191,
            d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207,
            d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223,
            d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239,
            d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255: in std_logic;
            S: in std_logic_vector (7 downto 0);
            r: out std_logic
        );
    end component;

    begin
        Mux256a1_0: Mux256a1 port map (d0(0), d1(0), d2(0), d3(0), d4(0), d5(0), d6(0), d7(0),
            d8(0), d9(0), d10(0), d11(0), d12(0), d13(0), d14(0), d15(0),
            d16(0), d17(0), d18(0), d19(0), d20(0), d21(0), d22(0), d23(0),
            d24(0), d25(0), d26(0), d27(0), d28(0), d29(0), d30(0), d31(0),
            d32(0), d33(0), d34(0), d35(0), d36(0), d37(0), d38(0), d39(0),
            d40(0), d41(0), d42(0), d43(0), d44(0), d45(0), d46(0), d47(0),
            d48(0), d49(0), d50(0), d51(0), d52(0), d53(0), d54(0), d55(0),
            d56(0), d57(0), d58(0), d59(0), d60(0), d61(0), d62(0), d63(0),
            d64(0), d65(0), d66(0), d67(0), d68(0), d69(0), d70(0), d71(0),
            d72(0), d73(0), d74(0), d75(0), d76(0), d77(0), d78(0), d79(0),
            d80(0), d81(0), d82(0), d83(0), d84(0), d85(0), d86(0), d87(0),
            d88(0), d89(0), d90(0), d91(0), d92(0), d93(0), d94(0), d95(0),
            d96(0), d97(0), d98(0), d99(0), d100(0), d101(0), d102(0), d103(0),
            d104(0), d105(0), d106(0), d107(0), d108(0), d109(0), d110(0), d111(0),
            d112(0), d113(0), d114(0), d115(0), d116(0), d117(0), d118(0), d119(0),
            d120(0), d121(0), d122(0), d123(0), d124(0), d125(0), d126(0), d127(0),
            d128(0), d129(0), d130(0), d131(0), d132(0), d133(0), d134(0), d135(0),
            d136(0), d137(0), d138(0), d139(0), d140(0), d141(0), d142(0), d143(0),
            d144(0), d145(0), d146(0), d147(0), d148(0), d149(0), d150(0), d151(0),
            d152(0), d153(0), d154(0), d155(0), d156(0), d157(0), d158(0), d159(0),
            d160(0), d161(0), d162(0), d163(0), d164(0), d165(0), d166(0), d167(0),
            d168(0), d169(0), d170(0), d171(0), d172(0), d173(0), d174(0), d175(0),
            d176(0), d177(0), d178(0), d179(0), d180(0), d181(0), d182(0), d183(0),
            d184(0), d185(0), d186(0), d187(0), d188(0), d189(0), d190(0), d191(0),
            d192(0), d193(0), d194(0), d195(0), d196(0), d197(0), d198(0), d199(0),
            d200(0), d201(0), d202(0), d203(0), d204(0), d205(0), d206(0), d207(0),
            d208(0), d209(0), d210(0), d211(0), d212(0), d213(0), d214(0), d215(0),
            d216(0), d217(0), d218(0), d219(0), d220(0), d221(0), d222(0), d223(0),
            d224(0), d225(0), d226(0), d227(0), d228(0), d229(0), d230(0), d231(0),
            d232(0), d233(0), d234(0), d235(0), d236(0), d237(0), d238(0), d239(0),
            d240(0), d241(0), d242(0), d243(0), d244(0), d245(0), d246(0), d247(0),
            d248(0), d249(0), d250(0), d251(0), d252(0), d253(0), d254(0), d255(0),
            S,
            r (0)
        );

        Mux256a1_1: Mux256a1 port map (d0(1), d1(1), d2(1), d3(1), d4(1), d5(1), d6(1), d7(1),
            d8(1), d9(1), d10(1), d11(1), d12(1), d13(1), d14(1), d15(1),
            d16(1), d17(1), d18(1), d19(1), d20(1), d21(1), d22(1), d23(1),
            d24(1), d25(1), d26(1), d27(1), d28(1), d29(1), d30(1), d31(1),
            d32(1), d33(1), d34(1), d35(1), d36(1), d37(1), d38(1), d39(1),
            d40(1), d41(1), d42(1), d43(1), d44(1), d45(1), d46(1), d47(1),
            d48(1), d49(1), d50(1), d51(1), d52(1), d53(1), d54(1), d55(1),
            d56(1), d57(1), d58(1), d59(1), d60(1), d61(1), d62(1), d63(1),
            d64(1), d65(1), d66(1), d67(1), d68(1), d69(1), d70(1), d71(1),
            d72(1), d73(1), d74(1), d75(1), d76(1), d77(1), d78(1), d79(1),
            d80(1), d81(1), d82(1), d83(1), d84(1), d85(1), d86(1), d87(1),
            d88(1), d89(1), d90(1), d91(1), d92(1), d93(1), d94(1), d95(1),
            d96(1), d97(1), d98(1), d99(1), d100(1), d101(1), d102(1), d103(1),
            d104(1), d105(1), d106(1), d107(1), d108(1), d109(1), d110(1), d111(1),
            d112(1), d113(1), d114(1), d115(1), d116(1), d117(1), d118(1), d119(1),
            d120(1), d121(1), d122(1), d123(1), d124(1), d125(1), d126(1), d127(1),
            d128(1), d129(1), d130(1), d131(1), d132(1), d133(1), d134(1), d135(1),
            d136(1), d137(1), d138(1), d139(1), d140(1), d141(1), d142(1), d143(1),
            d144(1), d145(1), d146(1), d147(1), d148(1), d149(1), d150(1), d151(1),
            d152(1), d153(1), d154(1), d155(1), d156(1), d157(1), d158(1), d159(1),
            d160(1), d161(1), d162(1), d163(1), d164(1), d165(1), d166(1), d167(1),
            d168(1), d169(1), d170(1), d171(1), d172(1), d173(1), d174(1), d175(1),
            d176(1), d177(1), d178(1), d179(1), d180(1), d181(1), d182(1), d183(1),
            d184(1), d185(1), d186(1), d187(1), d188(1), d189(1), d190(1), d191(1),
            d192(1), d193(1), d194(1), d195(1), d196(1), d197(1), d198(1), d199(1),
            d200(1), d201(1), d202(1), d203(1), d204(1), d205(1), d206(1), d207(1),
            d208(1), d209(1), d210(1), d211(1), d212(1), d213(1), d214(1), d215(1),
            d216(1), d217(1), d218(1), d219(1), d220(1), d221(1), d222(1), d223(1),
            d224(1), d225(1), d226(1), d227(1), d228(1), d229(1), d230(1), d231(1),
            d232(1), d233(1), d234(1), d235(1), d236(1), d237(1), d238(1), d239(1),
            d240(1), d241(1), d242(1), d243(1), d244(1), d245(1), d246(1), d247(1),
            d248(1), d249(1), d250(1), d251(1), d252(1), d253(1), d254(1), d255(1),
            S,
            r (1)
        );

        Mux256a1_2: Mux256a1 port map (d0(2), d1(2), d2(2), d3(2), d4(2), d5(2), d6(2), d7(2),
            d8(2), d9(2), d10(2), d11(2), d12(2), d13(2), d14(2), d15(2),
            d16(2), d17(2), d18(2), d19(2), d20(2), d21(2), d22(2), d23(2),
            d24(2), d25(2), d26(2), d27(2), d28(2), d29(2), d30(2), d31(2),
            d32(2), d33(2), d34(2), d35(2), d36(2), d37(2), d38(2), d39(2),
            d40(2), d41(2), d42(2), d43(2), d44(2), d45(2), d46(2), d47(2),
            d48(2), d49(2), d50(2), d51(2), d52(2), d53(2), d54(2), d55(2),
            d56(2), d57(2), d58(2), d59(2), d60(2), d61(2), d62(2), d63(2),
            d64(2), d65(2), d66(2), d67(2), d68(2), d69(2), d70(2), d71(2),
            d72(2), d73(2), d74(2), d75(2), d76(2), d77(2), d78(2), d79(2),
            d80(2), d81(2), d82(2), d83(2), d84(2), d85(2), d86(2), d87(2),
            d88(2), d89(2), d90(2), d91(2), d92(2), d93(2), d94(2), d95(2),
            d96(2), d97(2), d98(2), d99(2), d100(2), d101(2), d102(2), d103(2),
            d104(2), d105(2), d106(2), d107(2), d108(2), d109(2), d110(2), d111(2),
            d112(2), d113(2), d114(2), d115(2), d116(2), d117(2), d118(2), d119(2),
            d120(2), d121(2), d122(2), d123(2), d124(2), d125(2), d126(2), d127(2),
            d128(2), d129(2), d130(2), d131(2), d132(2), d133(2), d134(2), d135(2),
            d136(2), d137(2), d138(2), d139(2), d140(2), d141(2), d142(2), d143(2),
            d144(2), d145(2), d146(2), d147(2), d148(2), d149(2), d150(2), d151(2),
            d152(2), d153(2), d154(2), d155(2), d156(2), d157(2), d158(2), d159(2),
            d160(2), d161(2), d162(2), d163(2), d164(2), d165(2), d166(2), d167(2),
            d168(2), d169(2), d170(2), d171(2), d172(2), d173(2), d174(2), d175(2),
            d176(2), d177(2), d178(2), d179(2), d180(2), d181(2), d182(2), d183(2),
            d184(2), d185(2), d186(2), d187(2), d188(2), d189(2), d190(2), d191(2),
            d192(2), d193(2), d194(2), d195(2), d196(2), d197(2), d198(2), d199(2),
            d200(2), d201(2), d202(2), d203(2), d204(2), d205(2), d206(2), d207(2),
            d208(2), d209(2), d210(2), d211(2), d212(2), d213(2), d214(2), d215(2),
            d216(2), d217(2), d218(2), d219(2), d220(2), d221(2), d222(2), d223(2),
            d224(2), d225(2), d226(2), d227(2), d228(2), d229(2), d230(2), d231(2),
            d232(2), d233(2), d234(2), d235(2), d236(2), d237(2), d238(2), d239(2),
            d240(2), d241(2), d242(2), d243(2), d244(2), d245(2), d246(2), d247(2),
            d248(2), d249(2), d250(2), d251(2), d252(2), d253(2), d254(2), d255(2),
            S,
            r (2)
        );

        Mux256a1_3: Mux256a1 port map (d0(3), d1(3), d2(3), d3(3), d4(3), d5(3), d6(3), d7(3),
            d8(3), d9(3), d10(3), d11(3), d12(3), d13(3), d14(3), d15(3),
            d16(3), d17(3), d18(3), d19(3), d20(3), d21(3), d22(3), d23(3),
            d24(3), d25(3), d26(3), d27(3), d28(3), d29(3), d30(3), d31(3),
            d32(3), d33(3), d34(3), d35(3), d36(3), d37(3), d38(3), d39(3),
            d40(3), d41(3), d42(3), d43(3), d44(3), d45(3), d46(3), d47(3),
            d48(3), d49(3), d50(3), d51(3), d52(3), d53(3), d54(3), d55(3),
            d56(3), d57(3), d58(3), d59(3), d60(3), d61(3), d62(3), d63(3),
            d64(3), d65(3), d66(3), d67(3), d68(3), d69(3), d70(3), d71(3),
            d72(3), d73(3), d74(3), d75(3), d76(3), d77(3), d78(3), d79(3),
            d80(3), d81(3), d82(3), d83(3), d84(3), d85(3), d86(3), d87(3),
            d88(3), d89(3), d90(3), d91(3), d92(3), d93(3), d94(3), d95(3),
            d96(3), d97(3), d98(3), d99(3), d100(3), d101(3), d102(3), d103(3),
            d104(3), d105(3), d106(3), d107(3), d108(3), d109(3), d110(3), d111(3),
            d112(3), d113(3), d114(3), d115(3), d116(3), d117(3), d118(3), d119(3),
            d120(3), d121(3), d122(3), d123(3), d124(3), d125(3), d126(3), d127(3),
            d128(3), d129(3), d130(3), d131(3), d132(3), d133(3), d134(3), d135(3),
            d136(3), d137(3), d138(3), d139(3), d140(3), d141(3), d142(3), d143(3),
            d144(3), d145(3), d146(3), d147(3), d148(3), d149(3), d150(3), d151(3),
            d152(3), d153(3), d154(3), d155(3), d156(3), d157(3), d158(3), d159(3),
            d160(3), d161(3), d162(3), d163(3), d164(3), d165(3), d166(3), d167(3),
            d168(3), d169(3), d170(3), d171(3), d172(3), d173(3), d174(3), d175(3),
            d176(3), d177(3), d178(3), d179(3), d180(3), d181(3), d182(3), d183(3),
            d184(3), d185(3), d186(3), d187(3), d188(3), d189(3), d190(3), d191(3),
            d192(3), d193(3), d194(3), d195(3), d196(3), d197(3), d198(3), d199(3),
            d200(3), d201(3), d202(3), d203(3), d204(3), d205(3), d206(3), d207(3),
            d208(3), d209(3), d210(3), d211(3), d212(3), d213(3), d214(3), d215(3),
            d216(3), d217(3), d218(3), d219(3), d220(3), d221(3), d222(3), d223(3),
            d224(3), d225(3), d226(3), d227(3), d228(3), d229(3), d230(3), d231(3),
            d232(3), d233(3), d234(3), d235(3), d236(3), d237(3), d238(3), d239(3),
            d240(3), d241(3), d242(3), d243(3), d244(3), d245(3), d246(3), d247(3),
            d248(3), d249(3), d250(3), d251(3), d252(3), d253(3), d254(3), d255(3),
            S,
            r (3)
        );

        
        Mux256a1_4: Mux256a1 port map (d0(4), d1(4), d2(4), d3(4), d4(4), d5(4), d6(4), d7(4),
            d8(4), d9(4), d10(4), d11(4), d12(4), d13(4), d14(4), d15(4),
            d16(4), d17(4), d18(4), d19(4), d20(4), d21(4), d22(4), d23(4),
            d24(4), d25(4), d26(4), d27(4), d28(4), d29(4), d30(4), d31(4),
            d32(4), d33(4), d34(4), d35(4), d36(4), d37(4), d38(4), d39(4),
            d40(4), d41(4), d42(4), d43(4), d44(4), d45(4), d46(4), d47(4),
            d48(4), d49(4), d50(4), d51(4), d52(4), d53(4), d54(4), d55(4),
            d56(4), d57(4), d58(4), d59(4), d60(4), d61(4), d62(4), d63(4),
            d64(4), d65(4), d66(4), d67(4), d68(4), d69(4), d70(4), d71(4),
            d72(4), d73(4), d74(4), d75(4), d76(4), d77(4), d78(4), d79(4),
            d80(4), d81(4), d82(4), d83(4), d84(4), d85(4), d86(4), d87(4),
            d88(4), d89(4), d90(4), d91(4), d92(4), d93(4), d94(4), d95(4),
            d96(4), d97(4), d98(4), d99(4), d100(4), d101(4), d102(4), d103(4),
            d104(4), d105(4), d106(4), d107(4), d108(4), d109(4), d110(4), d111(4),
            d112(4), d113(4), d114(4), d115(4), d116(4), d117(4), d118(4), d119(4),
            d120(4), d121(4), d122(4), d123(4), d124(4), d125(4), d126(4), d127(4),
            d128(4), d129(4), d130(4), d131(4), d132(4), d133(4), d134(4), d135(4),
            d136(4), d137(4), d138(4), d139(4), d140(4), d141(4), d142(4), d143(4),
            d144(4), d145(4), d146(4), d147(4), d148(4), d149(4), d150(4), d151(4),
            d152(4), d153(4), d154(4), d155(4), d156(4), d157(4), d158(4), d159(4),
            d160(4), d161(4), d162(4), d163(4), d164(4), d165(4), d166(4), d167(4),
            d168(4), d169(4), d170(4), d171(4), d172(4), d173(4), d174(4), d175(4),
            d176(4), d177(4), d178(4), d179(4), d180(4), d181(4), d182(4), d183(4),
            d184(4), d185(4), d186(4), d187(4), d188(4), d189(4), d190(4), d191(4),
            d192(4), d193(4), d194(4), d195(4), d196(4), d197(4), d198(4), d199(4),
            d200(4), d201(4), d202(4), d203(4), d204(4), d205(4), d206(4), d207(4),
            d208(4), d209(4), d210(4), d211(4), d212(4), d213(4), d214(4), d215(4),
            d216(4), d217(4), d218(4), d219(4), d220(4), d221(4), d222(4), d223(4),
            d224(4), d225(4), d226(4), d227(4), d228(4), d229(4), d230(4), d231(4),
            d232(4), d233(4), d234(4), d235(4), d236(4), d237(4), d238(4), d239(4),
            d240(4), d241(4), d242(4), d243(4), d244(4), d245(4), d246(4), d247(4),
            d248(4), d249(4), d250(4), d251(4), d252(4), d253(4), d254(4), d255(4),
            S,
            r (4)
        );

        Mux256a1_5: Mux256a1 port map (d0(5), d1(5), d2(5), d3(5), d4(5), d5(5), d6(5), d7(5),
            d8(5), d9(5), d10(5), d11(5), d12(5), d13(5), d14(5), d15(5),
            d16(5), d17(5), d18(5), d19(5), d20(5), d21(5), d22(5), d23(5),
            d24(5), d25(5), d26(5), d27(5), d28(5), d29(5), d30(5), d31(5),
            d32(5), d33(5), d34(5), d35(5), d36(5), d37(5), d38(5), d39(5),
            d40(5), d41(5), d42(5), d43(5), d44(5), d45(5), d46(5), d47(5),
            d48(5), d49(5), d50(5), d51(5), d52(5), d53(5), d54(5), d55(5),
            d56(5), d57(5), d58(5), d59(5), d60(5), d61(5), d62(5), d63(5),
            d64(5), d65(5), d66(5), d67(5), d68(5), d69(5), d70(5), d71(5),
            d72(5), d73(5), d74(5), d75(5), d76(5), d77(5), d78(5), d79(5),
            d80(5), d81(5), d82(5), d83(5), d84(5), d85(5), d86(5), d87(5),
            d88(5), d89(5), d90(5), d91(5), d92(5), d93(5), d94(5), d95(5),
            d96(5), d97(5), d98(5), d99(5), d100(5), d101(5), d102(5), d103(5),
            d104(5), d105(5), d106(5), d107(5), d108(5), d109(5), d110(5), d111(5),
            d112(5), d113(5), d114(5), d115(5), d116(5), d117(5), d118(5), d119(5),
            d120(5), d121(5), d122(5), d123(5), d124(5), d125(5), d126(5), d127(5),
            d128(5), d129(5), d130(5), d131(5), d132(5), d133(5), d134(5), d135(5),
            d136(5), d137(5), d138(5), d139(5), d140(5), d141(5), d142(5), d143(5),
            d144(5), d145(5), d146(5), d147(5), d148(5), d149(5), d150(5), d151(5),
            d152(5), d153(5), d154(5), d155(5), d156(5), d157(5), d158(5), d159(5),
            d160(5), d161(5), d162(5), d163(5), d164(5), d165(5), d166(5), d167(5),
            d168(5), d169(5), d170(5), d171(5), d172(5), d173(5), d174(5), d175(5),
            d176(5), d177(5), d178(5), d179(5), d180(5), d181(5), d182(5), d183(5),
            d184(5), d185(5), d186(5), d187(5), d188(5), d189(5), d190(5), d191(5),
            d192(5), d193(5), d194(5), d195(5), d196(5), d197(5), d198(5), d199(5),
            d200(5), d201(5), d202(5), d203(5), d204(5), d205(5), d206(5), d207(5),
            d208(5), d209(5), d210(5), d211(5), d212(5), d213(5), d214(5), d215(5),
            d216(5), d217(5), d218(5), d219(5), d220(5), d221(5), d222(5), d223(5),
            d224(5), d225(5), d226(5), d227(5), d228(5), d229(5), d230(5), d231(5),
            d232(5), d233(5), d234(5), d235(5), d236(5), d237(5), d238(5), d239(5),
            d240(5), d241(5), d242(5), d243(5), d244(5), d245(5), d246(5), d247(5),
            d248(5), d249(5), d250(5), d251(5), d252(5), d253(5), d254(5), d255(5),
            S,
            r (5)
        );

        Mux256a1_6: Mux256a1 port map (d0(6), d1(6), d2(6), d3(6), d4(6), d5(6), d6(6), d7(6),
            d8(6), d9(6), d10(6), d11(6), d12(6), d13(6), d14(6), d15(6),
            d16(6), d17(6), d18(6), d19(6), d20(6), d21(6), d22(6), d23(6),
            d24(6), d25(6), d26(6), d27(6), d28(6), d29(6), d30(6), d31(6),
            d32(6), d33(6), d34(6), d35(6), d36(6), d37(6), d38(6), d39(6),
            d40(6), d41(6), d42(6), d43(6), d44(6), d45(6), d46(6), d47(6),
            d48(6), d49(6), d50(6), d51(6), d52(6), d53(6), d54(6), d55(6),
            d56(6), d57(6), d58(6), d59(6), d60(6), d61(6), d62(6), d63(6),
            d64(6), d65(6), d66(6), d67(6), d68(6), d69(6), d70(6), d71(6),
            d72(6), d73(6), d74(6), d75(6), d76(6), d77(6), d78(6), d79(6),
            d80(6), d81(6), d82(6), d83(6), d84(6), d85(6), d86(6), d87(6),
            d88(6), d89(6), d90(6), d91(6), d92(6), d93(6), d94(6), d95(6),
            d96(6), d97(6), d98(6), d99(6), d100(6), d101(6), d102(6), d103(6),
            d104(6), d105(6), d106(6), d107(6), d108(6), d109(6), d110(6), d111(6),
            d112(6), d113(6), d114(6), d115(6), d116(6), d117(6), d118(6), d119(6),
            d120(6), d121(6), d122(6), d123(6), d124(6), d125(6), d126(6), d127(6),
            d128(6), d129(6), d130(6), d131(6), d132(6), d133(6), d134(6), d135(6),
            d136(6), d137(6), d138(6), d139(6), d140(6), d141(6), d142(6), d143(6),
            d144(6), d145(6), d146(6), d147(6), d148(6), d149(6), d150(6), d151(6),
            d152(6), d153(6), d154(6), d155(6), d156(6), d157(6), d158(6), d159(6),
            d160(6), d161(6), d162(6), d163(6), d164(6), d165(6), d166(6), d167(6),
            d168(6), d169(6), d170(6), d171(6), d172(6), d173(6), d174(6), d175(6),
            d176(6), d177(6), d178(6), d179(6), d180(6), d181(6), d182(6), d183(6),
            d184(6), d185(6), d186(6), d187(6), d188(6), d189(6), d190(6), d191(6),
            d192(6), d193(6), d194(6), d195(6), d196(6), d197(6), d198(6), d199(6),
            d200(6), d201(6), d202(6), d203(6), d204(6), d205(6), d206(6), d207(6),
            d208(6), d209(6), d210(6), d211(6), d212(6), d213(6), d214(6), d215(6),
            d216(6), d217(6), d218(6), d219(6), d220(6), d221(6), d222(6), d223(6),
            d224(6), d225(6), d226(6), d227(6), d228(6), d229(6), d230(6), d231(6),
            d232(6), d233(6), d234(6), d235(6), d236(6), d237(6), d238(6), d239(6),
            d240(6), d241(6), d242(6), d243(6), d244(6), d245(6), d246(6), d247(6),
            d248(6), d249(6), d250(6), d251(6), d252(6), d253(6), d254(6), d255(6),
            S,
            r (6)
        );

        Mux256a1_7: Mux256a1 port map (d0(7), d1(7), d2(7), d3(7), d4(7), d5(7), d6(7), d7(7),
            d8(7), d9(7), d10(7), d11(7), d12(7), d13(7), d14(7), d15(7),
            d16(7), d17(7), d18(7), d19(7), d20(7), d21(7), d22(7), d23(7),
            d24(7), d25(7), d26(7), d27(7), d28(7), d29(7), d30(7), d31(7),
            d32(7), d33(7), d34(7), d35(7), d36(7), d37(7), d38(7), d39(7),
            d40(7), d41(7), d42(7), d43(7), d44(7), d45(7), d46(7), d47(7),
            d48(7), d49(7), d50(7), d51(7), d52(7), d53(7), d54(7), d55(7),
            d56(7), d57(7), d58(7), d59(7), d60(7), d61(7), d62(7), d63(7),
            d64(7), d65(7), d66(7), d67(7), d68(7), d69(7), d70(7), d71(7),
            d72(7), d73(7), d74(7), d75(7), d76(7), d77(7), d78(7), d79(7),
            d80(7), d81(7), d82(7), d83(7), d84(7), d85(7), d86(7), d87(7),
            d88(7), d89(7), d90(7), d91(7), d92(7), d93(7), d94(7), d95(7),
            d96(7), d97(7), d98(7), d99(7), d100(7), d101(7), d102(7), d103(7),
            d104(7), d105(7), d106(7), d107(7), d108(7), d109(7), d110(7), d111(7),
            d112(7), d113(7), d114(7), d115(7), d116(7), d117(7), d118(7), d119(7),
            d120(7), d121(7), d122(7), d123(7), d124(7), d125(7), d126(7), d127(7),
            d128(7), d129(7), d130(7), d131(7), d132(7), d133(7), d134(7), d135(7),
            d136(7), d137(7), d138(7), d139(7), d140(7), d141(7), d142(7), d143(7),
            d144(7), d145(7), d146(7), d147(7), d148(7), d149(7), d150(7), d151(7),
            d152(7), d153(7), d154(7), d155(7), d156(7), d157(7), d158(7), d159(7),
            d160(7), d161(7), d162(7), d163(7), d164(7), d165(7), d166(7), d167(7),
            d168(7), d169(7), d170(7), d171(7), d172(7), d173(7), d174(7), d175(7),
            d176(7), d177(7), d178(7), d179(7), d180(7), d181(7), d182(7), d183(7),
            d184(7), d185(7), d186(7), d187(7), d188(7), d189(7), d190(7), d191(7),
            d192(7), d193(7), d194(7), d195(7), d196(7), d197(7), d198(7), d199(7),
            d200(7), d201(7), d202(7), d203(7), d204(7), d205(7), d206(7), d207(7),
            d208(7), d209(7), d210(7), d211(7), d212(7), d213(7), d214(7), d215(7),
            d216(7), d217(7), d218(7), d219(7), d220(7), d221(7), d222(7), d223(7),
            d224(7), d225(7), d226(7), d227(7), d228(7), d229(7), d230(7), d231(7),
            d232(7), d233(7), d234(7), d235(7), d236(7), d237(7), d238(7), d239(7),
            d240(7), d241(7), d242(7), d243(7), d244(7), d245(7), d246(7), d247(7),
            d248(7), d249(7), d250(7), d251(7), d252(7), d253(7), d254(7), d255(7),
            S,
            r (7)
        );

        Mux256a1_8: Mux256a1 port map (
            d0(8), d1(8), d2(8), d3(8), d4(8), d5(8), d6(8), d7(8),
            d8(8), d9(8), d10(8), d11(8), d12(8), d13(8), d14(8), d15(8),
            d16(8), d17(8), d18(8), d19(8), d20(8), d21(8), d22(8), d23(8),
            d24(8), d25(8), d26(8), d27(8), d28(8), d29(8), d30(8), d31(8),
            d32(8), d33(8), d34(8), d35(8), d36(8), d37(8), d38(8), d39(8),
            d40(8), d41(8), d42(8), d43(8), d44(8), d45(8), d46(8), d47(8),
            d48(8), d49(8), d50(8), d51(8), d52(8), d53(8), d54(8), d55(8),
            d56(8), d57(8), d58(8), d59(8), d60(8), d61(8), d62(8), d63(8),
            d64(8), d65(8), d66(8), d67(8), d68(8), d69(8), d70(8), d71(8),
            d72(8), d73(8), d74(8), d75(8), d76(8), d77(8), d78(8), d79(8),
            d80(8), d81(8), d82(8), d83(8), d84(8), d85(8), d86(8), d87(8),
            d88(8), d89(8), d90(8), d91(8), d92(8), d93(8), d94(8), d95(8),
            d96(8), d97(8), d98(8), d99(8), d100(8), d101(8), d102(8), d103(8),
            d104(8), d105(8), d106(8), d107(8), d108(8), d109(8), d110(8), d111(8),
            d112(8), d113(8), d114(8), d115(8), d116(8), d117(8), d118(8), d119(8),
            d120(8), d121(8), d122(8), d123(8), d124(8), d125(8), d126(8), d127(8),
            d128(8), d129(8), d130(8), d131(8), d132(8), d133(8), d134(8), d135(8),
            d136(8), d137(8), d138(8), d139(8), d140(8), d141(8), d142(8), d143(8),
            d144(8), d145(8), d146(8), d147(8), d148(8), d149(8), d150(8), d151(8),
            d152(8), d153(8), d154(8), d155(8), d156(8), d157(8), d158(8), d159(8),
            d160(8), d161(8), d162(8), d163(8), d164(8), d165(8), d166(8), d167(8),
            d168(8), d169(8), d170(8), d171(8), d172(8), d173(8), d174(8), d175(8),
            d176(8), d177(8), d178(8), d179(8), d180(8), d181(8), d182(8), d183(8),
            d184(8), d185(8), d186(8), d187(8), d188(8), d189(8), d190(8), d191(8),
            d192(8), d193(8), d194(8), d195(8), d196(8), d197(8), d198(8), d199(8),
            d200(8), d201(8), d202(8), d203(8), d204(8), d205(8), d206(8), d207(8),
            d208(8), d209(8), d210(8), d211(8), d212(8), d213(8), d214(8), d215(8),
            d216(8), d217(8), d218(8), d219(8), d220(8), d221(8), d222(8), d223(8),
            d224(8), d225(8), d226(8), d227(8), d228(8), d229(8), d230(8), d231(8),
            d232(8), d233(8), d234(8), d235(8), d236(8), d237(8), d238(8), d239(8),
            d240(8), d241(8), d242(8), d243(8), d244(8), d245(8), d246(8), d247(8),
            d248(8), d249(8), d250(8), d251(8), d252(8), d253(8), d254(8), d255(8),
            S,
            r(8)
        );

        Mux256a1_9: Mux256a1 port map (
            d0(9), d1(9), d2(9), d3(9), d4(9), d5(9), d6(9), d7(9),
            d8(9), d9(9), d10(9), d11(9), d12(9), d13(9), d14(9), d15(9),
            d16(9), d17(9), d18(9), d19(9), d20(9), d21(9), d22(9), d23(9),
            d24(9), d25(9), d26(9), d27(9), d28(9), d29(9), d30(9), d31(9),
            d32(9), d33(9), d34(9), d35(9), d36(9), d37(9), d38(9), d39(9),
            d40(9), d41(9), d42(9), d43(9), d44(9), d45(9), d46(9), d47(9),
            d48(9), d49(9), d50(9), d51(9), d52(9), d53(9), d54(9), d55(9),
            d56(9), d57(9), d58(9), d59(9), d60(9), d61(9), d62(9), d63(9),
            d64(9), d65(9), d66(9), d67(9), d68(9), d69(9), d70(9), d71(9),
            d72(9), d73(9), d74(9), d75(9), d76(9), d77(9), d78(9), d79(9),
            d80(9), d81(9), d82(9), d83(9), d84(9), d85(9), d86(9), d87(9),
            d88(9), d89(9), d90(9), d91(9), d92(9), d93(9), d94(9), d95(9),
            d96(9), d97(9), d98(9), d99(9), d100(9), d101(9), d102(9), d103(9),
            d104(9), d105(9), d106(9), d107(9), d108(9), d109(9), d110(9), d111(9),
            d112(9), d113(9), d114(9), d115(9), d116(9), d117(9), d118(9), d119(9),
            d120(9), d121(9), d122(9), d123(9), d124(9), d125(9), d126(9), d127(9),
            d128(9), d129(9), d130(9), d131(9), d132(9), d133(9), d134(9), d135(9),
            d136(9), d137(9), d138(9), d139(9), d140(9), d141(9), d142(9), d143(9),
            d144(9), d145(9), d146(9), d147(9), d148(9), d149(9), d150(9), d151(9),
            d152(9), d153(9), d154(9), d155(9), d156(9), d157(9), d158(9), d159(9),
            d160(9), d161(9), d162(9), d163(9), d164(9), d165(9), d166(9), d167(9),
            d168(9), d169(9), d170(9), d171(9), d172(9), d173(9), d174(9), d175(9),
            d176(9), d177(9), d178(9), d179(9), d180(9), d181(9), d182(9), d183(9),
            d184(9), d185(9), d186(9), d187(9), d188(9), d189(9), d190(9), d191(9),
            d192(9), d193(9), d194(9), d195(9), d196(9), d197(9), d198(9), d199(9),
            d200(9), d201(9), d202(9), d203(9), d204(9), d205(9), d206(9), d207(9),
            d208(9), d209(9), d210(9), d211(9), d212(9), d213(9), d214(9), d215(9),
            d216(9), d217(9), d218(9), d219(9), d220(9), d221(9), d222(9), d223(9),
            d224(9), d225(9), d226(9), d227(9), d228(9), d229(9), d230(9), d231(9),
            d232(9), d233(9), d234(9), d235(9), d236(9), d237(9), d238(9), d239(9),
            d240(9), d241(9), d242(9), d243(9), d244(9), d245(9), d246(9), d247(9),
            d248(9), d249(9), d250(9), d251(9), d252(9), d253(9), d254(9), d255(9),
            S,
            r(9)
        );

        Mux256a1_10: Mux256a1 port map (
            d0(10), d1(10), d2(10), d3(10), d4(10), d5(10), d6(10), d7(10),
            d8(10), d9(10), d10(10), d11(10), d12(10), d13(10), d14(10), d15(10),
            d16(10), d17(10), d18(10), d19(10), d20(10), d21(10), d22(10), d23(10),
            d24(10), d25(10), d26(10), d27(10), d28(10), d29(10), d30(10), d31(10),
            d32(10), d33(10), d34(10), d35(10), d36(10), d37(10), d38(10), d39(10),
            d40(10), d41(10), d42(10), d43(10), d44(10), d45(10), d46(10), d47(10),
            d48(10), d49(10), d50(10), d51(10), d52(10), d53(10), d54(10), d55(10),
            d56(10), d57(10), d58(10), d59(10), d60(10), d61(10), d62(10), d63(10),
            d64(10), d65(10), d66(10), d67(10), d68(10), d69(10), d70(10), d71(10),
            d72(10), d73(10), d74(10), d75(10), d76(10), d77(10), d78(10), d79(10),
            d80(10), d81(10), d82(10), d83(10), d84(10), d85(10), d86(10), d87(10),
            d88(10), d89(10), d90(10), d91(10), d92(10), d93(10), d94(10), d95(10),
            d96(10), d97(10), d98(10), d99(10), d100(10), d101(10), d102(10), d103(10),
            d104(10), d105(10), d106(10), d107(10), d108(10), d109(10), d110(10), d111(10),
            d112(10), d113(10), d114(10), d115(10), d116(10), d117(10), d118(10), d119(10),
            d120(10), d121(10), d122(10), d123(10), d124(10), d125(10), d126(10), d127(10),
            d128(10), d129(10), d130(10), d131(10), d132(10), d133(10), d134(10), d135(10),
            d136(10), d137(10), d138(10), d139(10), d140(10), d141(10), d142(10), d143(10),
            d144(10), d145(10), d146(10), d147(10), d148(10), d149(10), d150(10), d151(10),
            d152(10), d153(10), d154(10), d155(10), d156(10), d157(10), d158(10), d159(10),
            d160(10), d161(10), d162(10), d163(10), d164(10), d165(10), d166(10), d167(10),
            d168(10), d169(10), d170(10), d171(10), d172(10), d173(10), d174(10), d175(10),
            d176(10), d177(10), d178(10), d179(10), d180(10), d181(10), d182(10), d183(10),
            d184(10), d185(10), d186(10), d187(10), d188(10), d189(10), d190(10), d191(10),
            d192(10), d193(10), d194(10), d195(10), d196(10), d197(10), d198(10), d199(10),
            d200(10), d201(10), d202(10), d203(10), d204(10), d205(10), d206(10), d207(10),
            d208(10), d209(10), d210(10), d211(10), d212(10), d213(10), d214(10), d215(10),
            d216(10), d217(10), d218(10), d219(10), d220(10), d221(10), d222(10), d223(10),
            d224(10), d225(10), d226(10), d227(10), d228(10), d229(10), d230(10), d231(10),
            d232(10), d233(10), d234(10), d235(10), d236(10), d237(10), d238(10), d239(10),
            d240(10), d241(10), d242(10), d243(10), d244(10), d245(10), d246(10), d247(10),
            d248(10), d249(10), d250(10), d251(10), d252(10), d253(10), d254(10), d255(10),
            S,
            r(10)
        );

        Mux256a1_11: Mux256a1 port map (
            d0(11), d1(11), d2(11), d3(11), d4(11), d5(11), d6(11), d7(11),
            d8(11), d9(11), d10(11), d11(11), d12(11), d13(11), d14(11), d15(11),
            d16(11), d17(11), d18(11), d19(11), d20(11), d21(11), d22(11), d23(11),
            d24(11), d25(11), d26(11), d27(11), d28(11), d29(11), d30(11), d31(11),
            d32(11), d33(11), d34(11), d35(11), d36(11), d37(11), d38(11), d39(11),
            d40(11), d41(11), d42(11), d43(11), d44(11), d45(11), d46(11), d47(11),
            d48(11), d49(11), d50(11), d51(11), d52(11), d53(11), d54(11), d55(11),
            d56(11), d57(11), d58(11), d59(11), d60(11), d61(11), d62(11), d63(11),
            d64(11), d65(11), d66(11), d67(11), d68(11), d69(11), d70(11), d71(11),
            d72(11), d73(11), d74(11), d75(11), d76(11), d77(11), d78(11), d79(11),
            d80(11), d81(11), d82(11), d83(11), d84(11), d85(11), d86(11), d87(11),
            d88(11), d89(11), d90(11), d91(11), d92(11), d93(11), d94(11), d95(11),
            d96(11), d97(11), d98(11), d99(11), d100(11), d101(11), d102(11), d103(11),
            d104(11), d105(11), d106(11), d107(11), d108(11), d109(11), d110(11), d111(11),
            d112(11), d113(11), d114(11), d115(11), d116(11), d117(11), d118(11), d119(11),
            d120(11), d121(11), d122(11), d123(11), d124(11), d125(11), d126(11), d127(11),
            d128(11), d129(11), d130(11), d131(11), d132(11), d133(11), d134(11), d135(11),
            d136(11), d137(11), d138(11), d139(11), d140(11), d141(11), d142(11), d143(11),
            d144(11), d145(11), d146(11), d147(11), d148(11), d149(11), d150(11), d151(11),
            d152(11), d153(11), d154(11), d155(11), d156(11), d157(11), d158(11), d159(11),
            d160(11), d161(11), d162(11), d163(11), d164(11), d165(11), d166(11), d167(11),
            d168(11), d169(11), d170(11), d171(11), d172(11), d173(11), d174(11), d175(11),
            d176(11), d177(11), d178(11), d179(11), d180(11), d181(11), d182(11), d183(11),
            d184(11), d185(11), d186(11), d187(11), d188(11), d189(11), d190(11), d191(11),
            d192(11), d193(11), d194(11), d195(11), d196(11), d197(11), d198(11), d199(11),
            d200(11), d201(11), d202(11), d203(11), d204(11), d205(11), d206(11), d207(11),
            d208(11), d209(11), d210(11), d211(11), d212(11), d213(11), d214(11), d215(11),
            d216(11), d217(11), d218(11), d219(11), d220(11), d221(11), d222(11), d223(11),
            d224(11), d225(11), d226(11), d227(11), d228(11), d229(11), d230(11), d231(11),
            d232(11), d233(11), d234(11), d235(11), d236(11), d237(11), d238(11), d239(11),
            d240(11), d241(11), d242(11), d243(11), d244(11), d245(11), d246(11), d247(11),
            d248(11), d249(11), d250(11), d251(11), d252(11), d253(11), d254(11), d255(11),
            S,
            r(11)
        );

        Mux256a1_12: Mux256a1 port map (
            d0(12), d1(12), d2(12), d3(12), d4(12), d5(12), d6(12), d7(12),
            d8(12), d9(12), d10(12), d11(12), d12(12), d13(12), d14(12), d15(12),
            d16(12), d17(12), d18(12), d19(12), d20(12), d21(12), d22(12), d23(12),
            d24(12), d25(12), d26(12), d27(12), d28(12), d29(12), d30(12), d31(12),
            d32(12), d33(12), d34(12), d35(12), d36(12), d37(12), d38(12), d39(12),
            d40(12), d41(12), d42(12), d43(12), d44(12), d45(12), d46(12), d47(12),
            d48(12), d49(12), d50(12), d51(12), d52(12), d53(12), d54(12), d55(12),
            d56(12), d57(12), d58(12), d59(12), d60(12), d61(12), d62(12), d63(12),
            d64(12), d65(12), d66(12), d67(12), d68(12), d69(12), d70(12), d71(12),
            d72(12), d73(12), d74(12), d75(12), d76(12), d77(12), d78(12), d79(12),
            d80(12), d81(12), d82(12), d83(12), d84(12), d85(12), d86(12), d87(12),
            d88(12), d89(12), d90(12), d91(12), d92(12), d93(12), d94(12), d95(12),
            d96(12), d97(12), d98(12), d99(12), d100(12), d101(12), d102(12), d103(12),
            d104(12), d105(12), d106(12), d107(12), d108(12), d109(12), d110(12), d111(12),
            d112(12), d113(12), d114(12), d115(12), d116(12), d117(12), d118(12), d119(12),
            d120(12), d121(12), d122(12), d123(12), d124(12), d125(12), d126(12), d127(12),
            d128(12), d129(12), d130(12), d131(12), d132(12), d133(12), d134(12), d135(12),
            d136(12), d137(12), d138(12), d139(12), d140(12), d141(12), d142(12), d143(12),
            d144(12), d145(12), d146(12), d147(12), d148(12), d149(12), d150(12), d151(12),
            d152(12), d153(12), d154(12), d155(12), d156(12), d157(12), d158(12), d159(12),
            d160(12), d161(12), d162(12), d163(12), d164(12), d165(12), d166(12), d167(12),
            d168(12), d169(12), d170(12), d171(12), d172(12), d173(12), d174(12), d175(12),
            d176(12), d177(12), d178(12), d179(12), d180(12), d181(12), d182(12), d183(12),
            d184(12), d185(12), d186(12), d187(12), d188(12), d189(12), d190(12), d191(12),
            d192(12), d193(12), d194(12), d195(12), d196(12), d197(12), d198(12), d199(12),
            d200(12), d201(12), d202(12), d203(12), d204(12), d205(12), d206(12), d207(12),
            d208(12), d209(12), d210(12), d211(12), d212(12), d213(12), d214(12), d215(12),
            d216(12), d217(12), d218(12), d219(12), d220(12), d221(12), d222(12), d223(12),
            d224(12), d225(12), d226(12), d227(12), d228(12), d229(12), d230(12), d231(12),
            d232(12), d233(12), d234(12), d235(12), d236(12), d237(12), d238(12), d239(12),
            d240(12), d241(12), d242(12), d243(12), d244(12), d245(12), d246(12), d247(12),
            d248(12), d249(12), d250(12), d251(12), d252(12), d253(12), d254(12), d255(12),
            S,
            r(12)
        );

        Mux256a1_13: Mux256a1 port map (
            d0(13), d1(13), d2(13), d3(13), d4(13), d5(13), d6(13), d7(13),
            d8(13), d9(13), d10(13), d11(13), d12(13), d13(13), d14(13), d15(13),
            d16(13), d17(13), d18(13), d19(13), d20(13), d21(13), d22(13), d23(13),
            d24(13), d25(13), d26(13), d27(13), d28(13), d29(13), d30(13), d31(13),
            d32(13), d33(13), d34(13), d35(13), d36(13), d37(13), d38(13), d39(13),
            d40(13), d41(13), d42(13), d43(13), d44(13), d45(13), d46(13), d47(13),
            d48(13), d49(13), d50(13), d51(13), d52(13), d53(13), d54(13), d55(13),
            d56(13), d57(13), d58(13), d59(13), d60(13), d61(13), d62(13), d63(13),
            d64(13), d65(13), d66(13), d67(13), d68(13), d69(13), d70(13), d71(13),
            d72(13), d73(13), d74(13), d75(13), d76(13), d77(13), d78(13), d79(13),
            d80(13), d81(13), d82(13), d83(13), d84(13), d85(13), d86(13), d87(13),
            d88(13), d89(13), d90(13), d91(13), d92(13), d93(13), d94(13), d95(13),
            d96(13), d97(13), d98(13), d99(13), d100(13), d101(13), d102(13), d103(13),
            d104(13), d105(13), d106(13), d107(13), d108(13), d109(13), d110(13), d111(13),
            d112(13), d113(13), d114(13), d115(13), d116(13), d117(13), d118(13), d119(13),
            d120(13), d121(13), d122(13), d123(13), d124(13), d125(13), d126(13), d127(13),
            d128(13), d129(13), d130(13), d131(13), d132(13), d133(13), d134(13), d135(13),
            d136(13), d137(13), d138(13), d139(13), d140(13), d141(13), d142(13), d143(13),
            d144(13), d145(13), d146(13), d147(13), d148(13), d149(13), d150(13), d151(13),
            d152(13), d153(13), d154(13), d155(13), d156(13), d157(13), d158(13), d159(13),
            d160(13), d161(13), d162(13), d163(13), d164(13), d165(13), d166(13), d167(13),
            d168(13), d169(13), d170(13), d171(13), d172(13), d173(13), d174(13), d175(13),
            d176(13), d177(13), d178(13), d179(13), d180(13), d181(13), d182(13), d183(13),
            d184(13), d185(13), d186(13), d187(13), d188(13), d189(13), d190(13), d191(13),
            d192(13), d193(13), d194(13), d195(13), d196(13), d197(13), d198(13), d199(13),
            d200(13), d201(13), d202(13), d203(13), d204(13), d205(13), d206(13), d207(13),
            d208(13), d209(13), d210(13), d211(13), d212(13), d213(13), d214(13), d215(13),
            d216(13), d217(13), d218(13), d219(13), d220(13), d221(13), d222(13), d223(13),
            d224(13), d225(13), d226(13), d227(13), d228(13), d229(13), d230(13), d231(13),
            d232(13), d233(13), d234(13), d235(13), d236(13), d237(13), d238(13), d239(13),
            d240(13), d241(13), d242(13), d243(13), d244(13), d245(13), d246(13), d247(13),
            d248(13), d249(13), d250(13), d251(13), d252(13), d253(13), d254(13), d255(13),
            S,
            r(13)
        );

        Mux256a1_14: Mux256a1 port map (
            d0(14), d1(14), d2(14), d3(14), d4(14), d5(14), d6(14), d7(14),
            d8(14), d9(14), d10(14), d11(14), d12(14), d13(14), d14(14), d15(14),
            d16(14), d17(14), d18(14), d19(14), d20(14), d21(14), d22(14), d23(14),
            d24(14), d25(14), d26(14), d27(14), d28(14), d29(14), d30(14), d31(14),
            d32(14), d33(14), d34(14), d35(14), d36(14), d37(14), d38(14), d39(14),
            d40(14), d41(14), d42(14), d43(14), d44(14), d45(14), d46(14), d47(14),
            d48(14), d49(14), d50(14), d51(14), d52(14), d53(14), d54(14), d55(14),
            d56(14), d57(14), d58(14), d59(14), d60(14), d61(14), d62(14), d63(14),
            d64(14), d65(14), d66(14), d67(14), d68(14), d69(14), d70(14), d71(14),
            d72(14), d73(14), d74(14), d75(14), d76(14), d77(14), d78(14), d79(14),
            d80(14), d81(14), d82(14), d83(14), d84(14), d85(14), d86(14), d87(14),
            d88(14), d89(14), d90(14), d91(14), d92(14), d93(14), d94(14), d95(14),
            d96(14), d97(14), d98(14), d99(14), d100(14), d101(14), d102(14), d103(14),
            d104(14), d105(14), d106(14), d107(14), d108(14), d109(14), d110(14), d111(14),
            d112(14), d113(14), d114(14), d115(14), d116(14), d117(14), d118(14), d119(14),
            d120(14), d121(14), d122(14), d123(14), d124(14), d125(14), d126(14), d127(14),
            d128(14), d129(14), d130(14), d131(14), d132(14), d133(14), d134(14), d135(14),
            d136(14), d137(14), d138(14), d139(14), d140(14), d141(14), d142(14), d143(14),
            d144(14), d145(14), d146(14), d147(14), d148(14), d149(14), d150(14), d151(14),
            d152(14), d153(14), d154(14), d155(14), d156(14), d157(14), d158(14), d159(14),
            d160(14), d161(14), d162(14), d163(14), d164(14), d165(14), d166(14), d167(14),
            d168(14), d169(14), d170(14), d171(14), d172(14), d173(14), d174(14), d175(14),
            d176(14), d177(14), d178(14), d179(14), d180(14), d181(14), d182(14), d183(14),
            d184(14), d185(14), d186(14), d187(14), d188(14), d189(14), d190(14), d191(14),
            d192(14), d193(14), d194(14), d195(14), d196(14), d197(14), d198(14), d199(14),
            d200(14), d201(14), d202(14), d203(14), d204(14), d205(14), d206(14), d207(14),
            d208(14), d209(14), d210(14), d211(14), d212(14), d213(14), d214(14), d215(14),
            d216(14), d217(14), d218(14), d219(14), d220(14), d221(14), d222(14), d223(14),
            d224(14), d225(14), d226(14), d227(14), d228(14), d229(14), d230(14), d231(14),
            d232(14), d233(14), d234(14), d235(14), d236(14), d237(14), d238(14), d239(14),
            d240(14), d241(14), d242(14), d243(14), d244(14), d245(14), d246(14), d247(14),
            d248(14), d249(14), d250(14), d251(14), d252(14), d253(14), d254(14), d255(14),
            S,
            r(14)
        );

        Mux256a1_15: Mux256a1 port map (
            d0(15), d1(15), d2(15), d3(15), d4(15), d5(15), d6(15), d7(15),
            d8(15), d9(15), d10(15), d11(15), d12(15), d13(15), d14(15), d15(15),
            d16(15), d17(15), d18(15), d19(15), d20(15), d21(15), d22(15), d23(15),
            d24(15), d25(15), d26(15), d27(15), d28(15), d29(15), d30(15), d31(15),
            d32(15), d33(15), d34(15), d35(15), d36(15), d37(15), d38(15), d39(15),
            d40(15), d41(15), d42(15), d43(15), d44(15), d45(15), d46(15), d47(15),
            d48(15), d49(15), d50(15), d51(15), d52(15), d53(15), d54(15), d55(15),
            d56(15), d57(15), d58(15), d59(15), d60(15), d61(15), d62(15), d63(15),
            d64(15), d65(15), d66(15), d67(15), d68(15), d69(15), d70(15), d71(15),
            d72(15), d73(15), d74(15), d75(15), d76(15), d77(15), d78(15), d79(15),
            d80(15), d81(15), d82(15), d83(15), d84(15), d85(15), d86(15), d87(15),
            d88(15), d89(15), d90(15), d91(15), d92(15), d93(15), d94(15), d95(15),
            d96(15), d97(15), d98(15), d99(15), d100(15), d101(15), d102(15), d103(15),
            d104(15), d105(15), d106(15), d107(15), d108(15), d109(15), d110(15), d111(15),
            d112(15), d113(15), d114(15), d115(15), d116(15), d117(15), d118(15), d119(15),
            d120(15), d121(15), d122(15), d123(15), d124(15), d125(15), d126(15), d127(15),
            d128(15), d129(15), d130(15), d131(15), d132(15), d133(15), d134(15), d135(15),
            d136(15), d137(15), d138(15), d139(15), d140(15), d141(15), d142(15), d143(15),
            d144(15), d145(15), d146(15), d147(15), d148(15), d149(15), d150(15), d151(15),
            d152(15), d153(15), d154(15), d155(15), d156(15), d157(15), d158(15), d159(15),
            d160(15), d161(15), d162(15), d163(15), d164(15), d165(15), d166(15), d167(15),
            d168(15), d169(15), d170(15), d171(15), d172(15), d173(15), d174(15), d175(15),
            d176(15), d177(15), d178(15), d179(15), d180(15), d181(15), d182(15), d183(15),
            d184(15), d185(15), d186(15), d187(15), d188(15), d189(15), d190(15), d191(15),
            d192(15), d193(15), d194(15), d195(15), d196(15), d197(15), d198(15), d199(15),
            d200(15), d201(15), d202(15), d203(15), d204(15), d205(15), d206(15), d207(15),
            d208(15), d209(15), d210(15), d211(15), d212(15), d213(15), d214(15), d215(15),
            d216(15), d217(15), d218(15), d219(15), d220(15), d221(15), d222(15), d223(15),
            d224(15), d225(15), d226(15), d227(15), d228(15), d229(15), d230(15), d231(15),
            d232(15), d233(15), d234(15), d235(15), d236(15), d237(15), d238(15), d239(15),
            d240(15), d241(15), d242(15), d243(15), d244(15), d245(15), d246(15), d247(15),
            d248(15), d249(15), d250(15), d251(15), d252(15), d253(15), d254(15), d255(15),
            S,
            r(15)
        );

        Mux256a1_16: Mux256a1 port map (
            d0(16), d1(16), d2(16), d3(16), d4(16), d5(16), d6(16), d7(16),
            d8(16), d9(16), d10(16), d11(16), d12(16), d13(16), d14(16), d15(16),
            d16(16), d17(16), d18(16), d19(16), d20(16), d21(16), d22(16), d23(16),
            d24(16), d25(16), d26(16), d27(16), d28(16), d29(16), d30(16), d31(16),
            d32(16), d33(16), d34(16), d35(16), d36(16), d37(16), d38(16), d39(16),
            d40(16), d41(16), d42(16), d43(16), d44(16), d45(16), d46(16), d47(16),
            d48(16), d49(16), d50(16), d51(16), d52(16), d53(16), d54(16), d55(16),
            d56(16), d57(16), d58(16), d59(16), d60(16), d61(16), d62(16), d63(16),
            d64(16), d65(16), d66(16), d67(16), d68(16), d69(16), d70(16), d71(16),
            d72(16), d73(16), d74(16), d75(16), d76(16), d77(16), d78(16), d79(16),
            d80(16), d81(16), d82(16), d83(16), d84(16), d85(16), d86(16), d87(16),
            d88(16), d89(16), d90(16), d91(16), d92(16), d93(16), d94(16), d95(16),
            d96(16), d97(16), d98(16), d99(16), d100(16), d101(16), d102(16), d103(16),
            d104(16), d105(16), d106(16), d107(16), d108(16), d109(16), d110(16), d111(16),
            d112(16), d113(16), d114(16), d115(16), d116(16), d117(16), d118(16), d119(16),
            d120(16), d121(16), d122(16), d123(16), d124(16), d125(16), d126(16), d127(16),
            d128(16), d129(16), d130(16), d131(16), d132(16), d133(16), d134(16), d135(16),
            d136(16), d137(16), d138(16), d139(16), d140(16), d141(16), d142(16), d143(16),
            d144(16), d145(16), d146(16), d147(16), d148(16), d149(16), d150(16), d151(16),
            d152(16), d153(16), d154(16), d155(16), d156(16), d157(16), d158(16), d159(16),
            d160(16), d161(16), d162(16), d163(16), d164(16), d165(16), d166(16), d167(16),
            d168(16), d169(16), d170(16), d171(16), d172(16), d173(16), d174(16), d175(16),
            d176(16), d177(16), d178(16), d179(16), d180(16), d181(16), d182(16), d183(16),
            d184(16), d185(16), d186(16), d187(16), d188(16), d189(16), d190(16), d191(16),
            d192(16), d193(16), d194(16), d195(16), d196(16), d197(16), d198(16), d199(16),
            d200(16), d201(16), d202(16), d203(16), d204(16), d205(16), d206(16), d207(16),
            d208(16), d209(16), d210(16), d211(16), d212(16), d213(16), d214(16), d215(16),
            d216(16), d217(16), d218(16), d219(16), d220(16), d221(16), d222(16), d223(16),
            d224(16), d225(16), d226(16), d227(16), d228(16), d229(16), d230(16), d231(16),
            d232(16), d233(16), d234(16), d235(16), d236(16), d237(16), d238(16), d239(16),
            d240(16), d241(16), d242(16), d243(16), d244(16), d245(16), d246(16), d247(16),
            d248(16), d249(16), d250(16), d251(16), d252(16), d253(16), d254(16), d255(16),
            S,
            r(16)
        );

        Mux256a1_17: Mux256a1 port map (
            d0(17), d1(17), d2(17), d3(17), d4(17), d5(17), d6(17), d7(17),
            d8(17), d9(17), d10(17), d11(17), d12(17), d13(17), d14(17), d15(17),
            d16(17), d17(17), d18(17), d19(17), d20(17), d21(17), d22(17), d23(17),
            d24(17), d25(17), d26(17), d27(17), d28(17), d29(17), d30(17), d31(17),
            d32(17), d33(17), d34(17), d35(17), d36(17), d37(17), d38(17), d39(17),
            d40(17), d41(17), d42(17), d43(17), d44(17), d45(17), d46(17), d47(17),
            d48(17), d49(17), d50(17), d51(17), d52(17), d53(17), d54(17), d55(17),
            d56(17), d57(17), d58(17), d59(17), d60(17), d61(17), d62(17), d63(17),
            d64(17), d65(17), d66(17), d67(17), d68(17), d69(17), d70(17), d71(17),
            d72(17), d73(17), d74(17), d75(17), d76(17), d77(17), d78(17), d79(17),
            d80(17), d81(17), d82(17), d83(17), d84(17), d85(17), d86(17), d87(17),
            d88(17), d89(17), d90(17), d91(17), d92(17), d93(17), d94(17), d95(17),
            d96(17), d97(17), d98(17), d99(17), d100(17), d101(17), d102(17), d103(17),
            d104(17), d105(17), d106(17), d107(17), d108(17), d109(17), d110(17), d111(17),
            d112(17), d113(17), d114(17), d115(17), d116(17), d117(17), d118(17), d119(17),
            d120(17), d121(17), d122(17), d123(17), d124(17), d125(17), d126(17), d127(17),
            d128(17), d129(17), d130(17), d131(17), d132(17), d133(17), d134(17), d135(17),
            d136(17), d137(17), d138(17), d139(17), d140(17), d141(17), d142(17), d143(17),
            d144(17), d145(17), d146(17), d147(17), d148(17), d149(17), d150(17), d151(17),
            d152(17), d153(17), d154(17), d155(17), d156(17), d157(17), d158(17), d159(17),
            d160(17), d161(17), d162(17), d163(17), d164(17), d165(17), d166(17), d167(17),
            d168(17), d169(17), d170(17), d171(17), d172(17), d173(17), d174(17), d175(17),
            d176(17), d177(17), d178(17), d179(17), d180(17), d181(17), d182(17), d183(17),
            d184(17), d185(17), d186(17), d187(17), d188(17), d189(17), d190(17), d191(17),
            d192(17), d193(17), d194(17), d195(17), d196(17), d197(17), d198(17), d199(17),
            d200(17), d201(17), d202(17), d203(17), d204(17), d205(17), d206(17), d207(17),
            d208(17), d209(17), d210(17), d211(17), d212(17), d213(17), d214(17), d215(17),
            d216(17), d217(17), d218(17), d219(17), d220(17), d221(17), d222(17), d223(17),
            d224(17), d225(17), d226(17), d227(17), d228(17), d229(17), d230(17), d231(17),
            d232(17), d233(17), d234(17), d235(17), d236(17), d237(17), d238(17), d239(17),
            d240(17), d241(17), d242(17), d243(17), d244(17), d245(17), d246(17), d247(17),
            d248(17), d249(17), d250(17), d251(17), d252(17), d253(17), d254(17), d255(17),
            S,
            r(17)
        );

        Mux256a1_18: Mux256a1 port map (
            d0(18), d1(18), d2(18), d3(18), d4(18), d5(18), d6(18), d7(18),
            d8(18), d9(18), d10(18), d11(18), d12(18), d13(18), d14(18), d15(18),
            d16(18), d17(18), d18(18), d19(18), d20(18), d21(18), d22(18), d23(18),
            d24(18), d25(18), d26(18), d27(18), d28(18), d29(18), d30(18), d31(18),
            d32(18), d33(18), d34(18), d35(18), d36(18), d37(18), d38(18), d39(18),
            d40(18), d41(18), d42(18), d43(18), d44(18), d45(18), d46(18), d47(18),
            d48(18), d49(18), d50(18), d51(18), d52(18), d53(18), d54(18), d55(18),
            d56(18), d57(18), d58(18), d59(18), d60(18), d61(18), d62(18), d63(18),
            d64(18), d65(18), d66(18), d67(18), d68(18), d69(18), d70(18), d71(18),
            d72(18), d73(18), d74(18), d75(18), d76(18), d77(18), d78(18), d79(18),
            d80(18), d81(18), d82(18), d83(18), d84(18), d85(18), d86(18), d87(18),
            d88(18), d89(18), d90(18), d91(18), d92(18), d93(18), d94(18), d95(18),
            d96(18), d97(18), d98(18), d99(18), d100(18), d101(18), d102(18), d103(18),
            d104(18), d105(18), d106(18), d107(18), d108(18), d109(18), d110(18), d111(18),
            d112(18), d113(18), d114(18), d115(18), d116(18), d117(18), d118(18), d119(18),
            d120(18), d121(18), d122(18), d123(18), d124(18), d125(18), d126(18), d127(18),
            d128(18), d129(18), d130(18), d131(18), d132(18), d133(18), d134(18), d135(18),
            d136(18), d137(18), d138(18), d139(18), d140(18), d141(18), d142(18), d143(18),
            d144(18), d145(18), d146(18), d147(18), d148(18), d149(18), d150(18), d151(18),
            d152(18), d153(18), d154(18), d155(18), d156(18), d157(18), d158(18), d159(18),
            d160(18), d161(18), d162(18), d163(18), d164(18), d165(18), d166(18), d167(18),
            d168(18), d169(18), d170(18), d171(18), d172(18), d173(18), d174(18), d175(18),
            d176(18), d177(18), d178(18), d179(18), d180(18), d181(18), d182(18), d183(18),
            d184(18), d185(18), d186(18), d187(18), d188(18), d189(18), d190(18), d191(18),
            d192(18), d193(18), d194(18), d195(18), d196(18), d197(18), d198(18), d199(18),
            d200(18), d201(18), d202(18), d203(18), d204(18), d205(18), d206(18), d207(18),
            d208(18), d209(18), d210(18), d211(18), d212(18), d213(18), d214(18), d215(18),
            d216(18), d217(18), d218(18), d219(18), d220(18), d221(18), d222(18), d223(18),
            d224(18), d225(18), d226(18), d227(18), d228(18), d229(18), d230(18), d231(18),
            d232(18), d233(18), d234(18), d235(18), d236(18), d237(18), d238(18), d239(18),
            d240(18), d241(18), d242(18), d243(18), d244(18), d245(18), d246(18), d247(18),
            d248(18), d249(18), d250(18), d251(18), d252(18), d253(18), d254(18), d255(18),
            S,
            r(18)
        );

        Mux256a1_19: Mux256a1 port map (
            d0(19), d1(19), d2(19), d3(19), d4(19), d5(19), d6(19), d7(19),
            d8(19), d9(19), d10(19), d11(19), d12(19), d13(19), d14(19), d15(19),
            d16(19), d17(19), d18(19), d19(19), d20(19), d21(19), d22(19), d23(19),
            d24(19), d25(19), d26(19), d27(19), d28(19), d29(19), d30(19), d31(19),
            d32(19), d33(19), d34(19), d35(19), d36(19), d37(19), d38(19), d39(19),
            d40(19), d41(19), d42(19), d43(19), d44(19), d45(19), d46(19), d47(19),
            d48(19), d49(19), d50(19), d51(19), d52(19), d53(19), d54(19), d55(19),
            d56(19), d57(19), d58(19), d59(19), d60(19), d61(19), d62(19), d63(19),
            d64(19), d65(19), d66(19), d67(19), d68(19), d69(19), d70(19), d71(19),
            d72(19), d73(19), d74(19), d75(19), d76(19), d77(19), d78(19), d79(19),
            d80(19), d81(19), d82(19), d83(19), d84(19), d85(19), d86(19), d87(19),
            d88(19), d89(19), d90(19), d91(19), d92(19), d93(19), d94(19), d95(19),
            d96(19), d97(19), d98(19), d99(19), d100(19), d101(19), d102(19), d103(19),
            d104(19), d105(19), d106(19), d107(19), d108(19), d109(19), d110(19), d111(19),
            d112(19), d113(19), d114(19), d115(19), d116(19), d117(19), d118(19), d119(19),
            d120(19), d121(19), d122(19), d123(19), d124(19), d125(19), d126(19), d127(19),
            d128(19), d129(19), d130(19), d131(19), d132(19), d133(19), d134(19), d135(19),
            d136(19), d137(19), d138(19), d139(19), d140(19), d141(19), d142(19), d143(19),
            d144(19), d145(19), d146(19), d147(19), d148(19), d149(19), d150(19), d151(19),
            d152(19), d153(19), d154(19), d155(19), d156(19), d157(19), d158(19), d159(19),
            d160(19), d161(19), d162(19), d163(19), d164(19), d165(19), d166(19), d167(19),
            d168(19), d169(19), d170(19), d171(19), d172(19), d173(19), d174(19), d175(19),
            d176(19), d177(19), d178(19), d179(19), d180(19), d181(19), d182(19), d183(19),
            d184(19), d185(19), d186(19), d187(19), d188(19), d189(19), d190(19), d191(19),
            d192(19), d193(19), d194(19), d195(19), d196(19), d197(19), d198(19), d199(19),
            d200(19), d201(19), d202(19), d203(19), d204(19), d205(19), d206(19), d207(19),
            d208(19), d209(19), d210(19), d211(19), d212(19), d213(19), d214(19), d215(19),
            d216(19), d217(19), d218(19), d219(19), d220(19), d221(19), d222(19), d223(19),
            d224(19), d225(19), d226(19), d227(19), d228(19), d229(19), d230(19), d231(19),
            d232(19), d233(19), d234(19), d235(19), d236(19), d237(19), d238(19), d239(19),
            d240(19), d241(19), d242(19), d243(19), d244(19), d245(19), d246(19), d247(19),
            d248(19), d249(19), d250(19), d251(19), d252(19), d253(19), d254(19), d255(19),
            S,
            r(19)
        );

        Mux256a1_20: Mux256a1 port map (
            d0(20), d1(20), d2(20), d3(20), d4(20), d5(20), d6(20), d7(20),
            d8(20), d9(20), d10(20), d11(20), d12(20), d13(20), d14(20), d15(20),
            d16(20), d17(20), d18(20), d19(20), d20(20), d21(20), d22(20), d23(20),
            d24(20), d25(20), d26(20), d27(20), d28(20), d29(20), d30(20), d31(20),
            d32(20), d33(20), d34(20), d35(20), d36(20), d37(20), d38(20), d39(20),
            d40(20), d41(20), d42(20), d43(20), d44(20), d45(20), d46(20), d47(20),
            d48(20), d49(20), d50(20), d51(20), d52(20), d53(20), d54(20), d55(20),
            d56(20), d57(20), d58(20), d59(20), d60(20), d61(20), d62(20), d63(20),
            d64(20), d65(20), d66(20), d67(20), d68(20), d69(20), d70(20), d71(20),
            d72(20), d73(20), d74(20), d75(20), d76(20), d77(20), d78(20), d79(20),
            d80(20), d81(20), d82(20), d83(20), d84(20), d85(20), d86(20), d87(20),
            d88(20), d89(20), d90(20), d91(20), d92(20), d93(20), d94(20), d95(20),
            d96(20), d97(20), d98(20), d99(20), d100(20), d101(20), d102(20), d103(20),
            d104(20), d105(20), d106(20), d107(20), d108(20), d109(20), d110(20), d111(20),
            d112(20), d113(20), d114(20), d115(20), d116(20), d117(20), d118(20), d119(20),
            d120(20), d121(20), d122(20), d123(20), d124(20), d125(20), d126(20), d127(20),
            d128(20), d129(20), d130(20), d131(20), d132(20), d133(20), d134(20), d135(20),
            d136(20), d137(20), d138(20), d139(20), d140(20), d141(20), d142(20), d143(20),
            d144(20), d145(20), d146(20), d147(20), d148(20), d149(20), d150(20), d151(20),
            d152(20), d153(20), d154(20), d155(20), d156(20), d157(20), d158(20), d159(20),
            d160(20), d161(20), d162(20), d163(20), d164(20), d165(20), d166(20), d167(20),
            d168(20), d169(20), d170(20), d171(20), d172(20), d173(20), d174(20), d175(20),
            d176(20), d177(20), d178(20), d179(20), d180(20), d181(20), d182(20), d183(20),
            d184(20), d185(20), d186(20), d187(20), d188(20), d189(20), d190(20), d191(20),
            d192(20), d193(20), d194(20), d195(20), d196(20), d197(20), d198(20), d199(20),
            d200(20), d201(20), d202(20), d203(20), d204(20), d205(20), d206(20), d207(20),
            d208(20), d209(20), d210(20), d211(20), d212(20), d213(20), d214(20), d215(20),
            d216(20), d217(20), d218(20), d219(20), d220(20), d221(20), d222(20), d223(20),
            d224(20), d225(20), d226(20), d227(20), d228(20), d229(20), d230(20), d231(20),
            d232(20), d233(20), d234(20), d235(20), d236(20), d237(20), d238(20), d239(20),
            d240(20), d241(20), d242(20), d243(20), d244(20), d245(20), d246(20), d247(20),
            d248(20), d249(20), d250(20), d251(20), d252(20), d253(20), d254(20), d255(20),
            S,
            r(20)
        );

        Mux256a1_21: Mux256a1 port map (
            d0(21), d1(21), d2(21), d3(21), d4(21), d5(21), d6(21), d7(21),
            d8(21), d9(21), d10(21), d11(21), d12(21), d13(21), d14(21), d15(21),
            d16(21), d17(21), d18(21), d19(21), d20(21), d21(21), d22(21), d23(21),
            d24(21), d25(21), d26(21), d27(21), d28(21), d29(21), d30(21), d31(21),
            d32(21), d33(21), d34(21), d35(21), d36(21), d37(21), d38(21), d39(21),
            d40(21), d41(21), d42(21), d43(21), d44(21), d45(21), d46(21), d47(21),
            d48(21), d49(21), d50(21), d51(21), d52(21), d53(21), d54(21), d55(21),
            d56(21), d57(21), d58(21), d59(21), d60(21), d61(21), d62(21), d63(21),
            d64(21), d65(21), d66(21), d67(21), d68(21), d69(21), d70(21), d71(21),
            d72(21), d73(21), d74(21), d75(21), d76(21), d77(21), d78(21), d79(21),
            d80(21), d81(21), d82(21), d83(21), d84(21), d85(21), d86(21), d87(21),
            d88(21), d89(21), d90(21), d91(21), d92(21), d93(21), d94(21), d95(21),
            d96(21), d97(21), d98(21), d99(21), d100(21), d101(21), d102(21), d103(21),
            d104(21), d105(21), d106(21), d107(21), d108(21), d109(21), d110(21), d111(21),
            d112(21), d113(21), d114(21), d115(21), d116(21), d117(21), d118(21), d119(21),
            d120(21), d121(21), d122(21), d123(21), d124(21), d125(21), d126(21), d127(21),
            d128(21), d129(21), d130(21), d131(21), d132(21), d133(21), d134(21), d135(21),
            d136(21), d137(21), d138(21), d139(21), d140(21), d141(21), d142(21), d143(21),
            d144(21), d145(21), d146(21), d147(21), d148(21), d149(21), d150(21), d151(21),
            d152(21), d153(21), d154(21), d155(21), d156(21), d157(21), d158(21), d159(21),
            d160(21), d161(21), d162(21), d163(21), d164(21), d165(21), d166(21), d167(21),
            d168(21), d169(21), d170(21), d171(21), d172(21), d173(21), d174(21), d175(21),
            d176(21), d177(21), d178(21), d179(21), d180(21), d181(21), d182(21), d183(21),
            d184(21), d185(21), d186(21), d187(21), d188(21), d189(21), d190(21), d191(21),
            d192(21), d193(21), d194(21), d195(21), d196(21), d197(21), d198(21), d199(21),
            d200(21), d201(21), d202(21), d203(21), d204(21), d205(21), d206(21), d207(21),
            d208(21), d209(21), d210(21), d211(21), d212(21), d213(21), d214(21), d215(21),
            d216(21), d217(21), d218(21), d219(21), d220(21), d221(21), d222(21), d223(21),
            d224(21), d225(21), d226(21), d227(21), d228(21), d229(21), d230(21), d231(21),
            d232(21), d233(21), d234(21), d235(21), d236(21), d237(21), d238(21), d239(21),
            d240(21), d241(21), d242(21), d243(21), d244(21), d245(21), d246(21), d247(21),
            d248(21), d249(21), d250(21), d251(21), d252(21), d253(21), d254(21), d255(21),
            S,
            r(21)
        );

        Mux256a1_22: Mux256a1 port map (
            d0(22), d1(22), d2(22), d3(22), d4(22), d5(22), d6(22), d7(22),
            d8(22), d9(22), d10(22), d11(22), d12(22), d13(22), d14(22), d15(22),
            d16(22), d17(22), d18(22), d19(22), d20(22), d21(22), d22(22), d23(22),
            d24(22), d25(22), d26(22), d27(22), d28(22), d29(22), d30(22), d31(22),
            d32(22), d33(22), d34(22), d35(22), d36(22), d37(22), d38(22), d39(22),
            d40(22), d41(22), d42(22), d43(22), d44(22), d45(22), d46(22), d47(22),
            d48(22), d49(22), d50(22), d51(22), d52(22), d53(22), d54(22), d55(22),
            d56(22), d57(22), d58(22), d59(22), d60(22), d61(22), d62(22), d63(22),
            d64(22), d65(22), d66(22), d67(22), d68(22), d69(22), d70(22), d71(22),
            d72(22), d73(22), d74(22), d75(22), d76(22), d77(22), d78(22), d79(22),
            d80(22), d81(22), d82(22), d83(22), d84(22), d85(22), d86(22), d87(22),
            d88(22), d89(22), d90(22), d91(22), d92(22), d93(22), d94(22), d95(22),
            d96(22), d97(22), d98(22), d99(22), d100(22), d101(22), d102(22), d103(22),
            d104(22), d105(22), d106(22), d107(22), d108(22), d109(22), d110(22), d111(22),
            d112(22), d113(22), d114(22), d115(22), d116(22), d117(22), d118(22), d119(22),
            d120(22), d121(22), d122(22), d123(22), d124(22), d125(22), d126(22), d127(22),
            d128(22), d129(22), d130(22), d131(22), d132(22), d133(22), d134(22), d135(22),
            d136(22), d137(22), d138(22), d139(22), d140(22), d141(22), d142(22), d143(22),
            d144(22), d145(22), d146(22), d147(22), d148(22), d149(22), d150(22), d151(22),
            d152(22), d153(22), d154(22), d155(22), d156(22), d157(22), d158(22), d159(22),
            d160(22), d161(22), d162(22), d163(22), d164(22), d165(22), d166(22), d167(22),
            d168(22), d169(22), d170(22), d171(22), d172(22), d173(22), d174(22), d175(22),
            d176(22), d177(22), d178(22), d179(22), d180(22), d181(22), d182(22), d183(22),
            d184(22), d185(22), d186(22), d187(22), d188(22), d189(22), d190(22), d191(22),
            d192(22), d193(22), d194(22), d195(22), d196(22), d197(22), d198(22), d199(22),
            d200(22), d201(22), d202(22), d203(22), d204(22), d205(22), d206(22), d207(22),
            d208(22), d209(22), d210(22), d211(22), d212(22), d213(22), d214(22), d215(22),
            d216(22), d217(22), d218(22), d219(22), d220(22), d221(22), d222(22), d223(22),
            d224(22), d225(22), d226(22), d227(22), d228(22), d229(22), d230(22), d231(22),
            d232(22), d233(22), d234(22), d235(22), d236(22), d237(22), d238(22), d239(22),
            d240(22), d241(22), d242(22), d243(22), d244(22), d245(22), d246(22), d247(22),
            d248(22), d249(22), d250(22), d251(22), d252(22), d253(22), d254(22), d255(22),
            S,
            r(22)
        );

    Mux256a1_23: Mux256a1 port map (
        d0(23), d1(23), d2(23), d3(23), d4(23), d5(23), d6(23), d7(23),
        d8(23), d9(23), d10(23), d11(23), d12(23), d13(23), d14(23), d15(23),
        d16(23), d17(23), d18(23), d19(23), d20(23), d21(23), d22(23), d23(23),
        d24(23), d25(23), d26(23), d27(23), d28(23), d29(23), d30(23), d31(23),
        d32(23), d33(23), d34(23), d35(23), d36(23), d37(23), d38(23), d39(23),
        d40(23), d41(23), d42(23), d43(23), d44(23), d45(23), d46(23), d47(23),
        d48(23), d49(23), d50(23), d51(23), d52(23), d53(23), d54(23), d55(23),
        d56(23), d57(23), d58(23), d59(23), d60(23), d61(23), d62(23), d63(23),
        d64(23), d65(23), d66(23), d67(23), d68(23), d69(23), d70(23), d71(23),
        d72(23), d73(23), d74(23), d75(23), d76(23), d77(23), d78(23), d79(23),
        d80(23), d81(23), d82(23), d83(23), d84(23), d85(23), d86(23), d87(23),
        d88(23), d89(23), d90(23), d91(23), d92(23), d93(23), d94(23), d95(23),
        d96(23), d97(23), d98(23), d99(23), d100(23), d101(23), d102(23), d103(23),
        d104(23), d105(23), d106(23), d107(23), d108(23), d109(23), d110(23), d111(23),
        d112(23), d113(23), d114(23), d115(23), d116(23), d117(23), d118(23), d119(23),
        d120(23), d121(23), d122(23), d123(23), d124(23), d125(23), d126(23), d127(23),
        d128(23), d129(23), d130(23), d131(23), d132(23), d133(23), d134(23), d135(23),
        d136(23), d137(23), d138(23), d139(23), d140(23), d141(23), d142(23), d143(23),
        d144(23), d145(23), d146(23), d147(23), d148(23), d149(23), d150(23), d151(23),
        d152(23), d153(23), d154(23), d155(23), d156(23), d157(23), d158(23), d159(23),
        d160(23), d161(23), d162(23), d163(23), d164(23), d165(23), d166(23), d167(23),
        d168(23), d169(23), d170(23), d171(23), d172(23), d173(23), d174(23), d175(23),
        d176(23), d177(23), d178(23), d179(23), d180(23), d181(23), d182(23), d183(23),
        d184(23), d185(23), d186(23), d187(23), d188(23), d189(23), d190(23), d191(23),
        d192(23), d193(23), d194(23), d195(23), d196(23), d197(23), d198(23), d199(23),
        d200(23), d201(23), d202(23), d203(23), d204(23), d205(23), d206(23), d207(23),
        d208(23), d209(23), d210(23), d211(23), d212(23), d213(23), d214(23), d215(23),
        d216(23), d217(23), d218(23), d219(23), d220(23), d221(23), d222(23), d223(23),
        d224(23), d225(23), d226(23), d227(23), d228(23), d229(23), d230(23), d231(23),
        d232(23), d233(23), d234(23), d235(23), d236(23), d237(23), d238(23), d239(23),
        d240(23), d241(23), d242(23), d243(23), d244(23), d245(23), d246(23), d247(23),
        d248(23), d249(23), d250(23), d251(23), d252(23), d253(23), d254(23), d255(23),
        S,
        r(23)
    );


    Mux256a1_24: Mux256a1 port map (
        d0(24), d1(24), d2(24), d3(24), d4(24), d5(24), d6(24), d7(24),
        d8(24), d9(24), d10(24), d11(24), d12(24), d13(24), d14(24), d15(24),
        d16(24), d17(24), d18(24), d19(24), d20(24), d21(24), d22(24), d23(24),
        d24(24), d25(24), d26(24), d27(24), d28(24), d29(24), d30(24), d31(24),
        d32(24), d33(24), d34(24), d35(24), d36(24), d37(24), d38(24), d39(24),
        d40(24), d41(24), d42(24), d43(24), d44(24), d45(24), d46(24), d47(24),
        d48(24), d49(24), d50(24), d51(24), d52(24), d53(24), d54(24), d55(24),
        d56(24), d57(24), d58(24), d59(24), d60(24), d61(24), d62(24), d63(24),
        d64(24), d65(24), d66(24), d67(24), d68(24), d69(24), d70(24), d71(24),
        d72(24), d73(24), d74(24), d75(24), d76(24), d77(24), d78(24), d79(24),
        d80(24), d81(24), d82(24), d83(24), d84(24), d85(24), d86(24), d87(24),
        d88(24), d89(24), d90(24), d91(24), d92(24), d93(24), d94(24), d95(24),
        d96(24), d97(24), d98(24), d99(24), d100(24), d101(24), d102(24), d103(24),
        d104(24), d105(24), d106(24), d107(24), d108(24), d109(24), d110(24), d111(24),
        d112(24), d113(24), d114(24), d115(24), d116(24), d117(24), d118(24), d119(24),
        d120(24), d121(24), d122(24), d123(24), d124(24), d125(24), d126(24), d127(24),
        d128(24), d129(24), d130(24), d131(24), d132(24), d133(24), d134(24), d135(24),
        d136(24), d137(24), d138(24), d139(24), d140(24), d141(24), d142(24), d143(24),
        d144(24), d145(24), d146(24), d147(24), d148(24), d149(24), d150(24), d151(24),
        d152(24), d153(24), d154(24), d155(24), d156(24), d157(24), d158(24), d159(24),
        d160(24), d161(24), d162(24), d163(24), d164(24), d165(24), d166(24), d167(24),
        d168(24), d169(24), d170(24), d171(24), d172(24), d173(24), d174(24), d175(24),
        d176(24), d177(24), d178(24), d179(24), d180(24), d181(24), d182(24), d183(24),
        d184(24), d185(24), d186(24), d187(24), d188(24), d189(24), d190(24), d191(24),
        d192(24), d193(24), d194(24), d195(24), d196(24), d197(24), d198(24), d199(24),
        d200(24), d201(24), d202(24), d203(24), d204(24), d205(24), d206(24), d207(24),
        d208(24), d209(24), d210(24), d211(24), d212(24), d213(24), d214(24), d215(24),
        d216(24), d217(24), d218(24), d219(24), d220(24), d221(24), d222(24), d223(24),
        d224(24), d225(24), d226(24), d227(24), d228(24), d229(24), d230(24), d231(24),
        d232(24), d233(24), d234(24), d235(24), d236(24), d237(24), d238(24), d239(24),
        d240(24), d241(24), d242(24), d243(24), d244(24), d245(24), d246(24), d247(24),
        d248(24), d249(24), d250(24), d251(24), d252(24), d253(24), d254(24), d255(24),
        S,
        r(24)
    );





    end architecture;